��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���G�H�ƻ	�"�iQ�����3�7Q��㼫F|�ݽ0��@h ���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�s8�R�	�}����i�'������\�N
x��]Qu ������[���a�8%`��4�s�6�XAoeuxLZ�#8�d~O�GӔ�<4��ˌ�ň��h��=i�@x_\q�jB�Fg�Y씤`��p�܂aQ�"6�l�:��3�����U���T���딣0&_���X0���2|	p��rw@	@us���
���m�jm\J�ԭyq�`݊�|���"rG�
���}�\�.�DV	��dU�;�\�]���џ�_�v%�]��4�:j�l�,9��I{��8�H��s8[Z��pM�i?��n;�|-���g]�ܜ�׫��$R7�t��q�t,�,v*5���a["<7U�i�#!����P�>�>��2$u�{}�=�vsO�~�fB��z��35{���fqx>�a����FIҶn��JٕTm7�+���%U����Ǘ�Y�@�:t''�#w��E�N���q�pH��5�+F�DÀ��h�)4�B��ٴy�@�Wx+�-EP,]�!�`�(i3!�`�(i3�=��W@&��?N����������/�}���1�1�ҕ�/37���E�D��`X��$D@P�a;����XV��w�K�	�f<���V��m̖n�Uvsȸ�"rR!�`�(i3��6��*}���l4�$�(�����ȍW�j��RB��4���O�>�k}�r���ۑQEYx�q�;��{C��c�S+d�J�Г��f�u�����!-��B<ԧ�[��+��sȸ�"rR!�`�(i3�B�'��a�{�ç�o�����0����(R\֎u��� Sgȼ�sʫ|H�ͩ�QϿ�ey��<0!�`�(i3!�`�(i3����N����������(��K.�j��RB{?a� ~>>ը܅%Gbغ���:�9I�uEd�=�WT�%�i���*��W~�O�N����X����3�ok!�`�(i3!�`�(i3������!���C�/�y���ܴ�WM�P[��j�$�*7I���y�L�=sȸ�"rR!�`�(i3�2 /��u��
���ƸtU�����3�(�^��o�D24N<I8����\.Wֵ*&E�^8��xt��:_/�~8����A�߲wLB�w���#✲�@�킍�"�?���Fz�!�`�(i3!�`�(i3L�E��1I�OfUA`���B��ҙ����WH%���ܜ?n昼�2#:�^��R�8���2O��'HY-w�Y��k��ı����~K�%���c)�ӣ4��Ny5�7\F���r��RL�a)����c���,�%���pY�� e�o�"��Ը��w�>��S9�����}����j���k�8���҆�|n����:Vx�p*+i#GBp�K�K%��2��ѕ���^�4㥭����!�9�R��zF�YQ��s,�~TM�e�w�G��7�"���`�[����Y�1m���	�ۚ0������}n)�Z�:���*S9���ݬ�NY���eb��D@f$�Ƣ�/�?�� �@ǜ7�\3���8�{�0]�P:�Qu��w)�S-!�����c�J�M=�!FLL4��)(�"`z8�:r&@�G	���su�]bu̎x4�J����4�����
� �AH�*��.�/7� GD��O�etwa�¢>�P��ѕ���5��ˬ�d�>]@a��X��zorL�o5'�� ��,Iw�)������\�4�si�W���y(;⟝*#X{g�n}�y�mq��o?�M��;]�_8����@�r��_��{,!.��m�!=�y����h�}y(;⟝*#X{g�n}�y��i�]w�o?�M��;]ԙ���!�4<�`�H��B��͌�a^X����\�4�si�W���)���32*D�S�ar���!�@C�Sd,�ϱ��|�GJ Ւ�&��(\+�5e��q���H�!j�h_}�������5�6�tR��\�4�si�W���jh�6g�*D�S�ar!���1��Sd,�ϱ��N��[r�����M�jT��#�)��Q=����n*99�!/����RL�a)8��Q̮����i�P�u3 ����YZX��w�>��S�rA��0Ǧ,\ަ�It���[���*\��_���w﴾�J]�r4EG�j��f6&��?N����l	��n����j�t�A�-*�Y��
Ż�y�Qg>7��^�V�Ϟ��^�ڥ���a����iO��ޔUH�>�r�O��C��0����"'��/��I��$MAF�)�hg���!�zg�Z�$;���D��T���=c��D�P��S���D���i����	x]�<���e8ưc��L�F�f��ӕ� +u��IPu���V��XO�����y�k[��K;���\�4�sR���i1�8Y�&�\��\�õɆ#�Ԗ̋n;�q�m
cxFu�n����RF�g�ï;K6�{�jc�^�p����"��J�Zj����l�� q#��RL�a)8��Q̮��,�%��/w����M��oսw�>��SU��Pa����4#!(��*/�|�v������J��\���a6�Ͳ
�3�K,��,Iw�)�K�������	x]̍��;��8ưc�꿷i=��䏇W��s�!5�Edɲ�<a�l�y@���lk�߻�<��F[����N���5���ݱ�A�fܑלoJ|��\�4�s��{��]Q�TT	q��$��<�z5��J��eb�hW!'!7U�i�#!����P�>;�Ղ��G}Z��2�p��Oi�v���j�������JM�7")�E�'3H��[e)�p�R\��ꫜp&C����/B!,�G�;(�B�T0�z$�}���E6sC&�gG��Hc�e$���=M��8�w'��(�D�&�〨����cZ	�M2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vce��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc/?�s�m/C�Ѽ?��Q2�=W�֯�^��N�&��^˻f��	g�y���}�ZC��aNvA�;�m�\��qi��p�7���I�4�Ȧ5
�
Tt˩�e�J�4>��1lD�J8���=Udq��D��tw:g+��T��d^��_|��3g�ݜ��s8[Z�`
5��*�z�������D���J7"z��cX��aC�h�>�N{a�9Ow�Y��k��ı����~K�%���c)�ӣ4�"�却G�����d���q����c��� �7ht��}j"�,�>E��4];ˍH�!�`�(i3MP$���p�B��F��|��v�0<๸u�Ґ�eb�3���)�[���6JHn��z��x�f7﹏T?�7G|`}���@/��(�ߜ1��E����F�'n�^0o"�,�>E��� ����{7$0~'��&\VI`,�ʺ�;[��\�v�!�`�(i3p40�zɈ�Ќ��*��4.���Xt�.U��'n�^0o"�,�>E���$�F�s+���!,�U&��/�,�#�H�1c����O}����g�a!�`�(i3!�`�(i3!�`�(i3!�`�(i3<�6�Q=@^7&ģM:�5t�W?pk� �,�� �0r��*�'yV��>���_��l���׷fh����y����vG\��o�&��v�/��k�����.����$`0�S����[LKS}?���\z-ܘ�u}����зq8�ЈR���b�>��;C@������9qj�xm�N��p��ٸ�z��������� ͢��8k��T9s*ox!�Q�W��ݚ�Н�!�`�(i3!�`�(i3!�`�(i3!�`�(i3��7zgN<�|�taf��P���p�Y�Es�D��P+G2�9��?���\z-��EM���
+����r"�,�>E��4];ˍH�!�`�(i3��y�s���	L'J����Rb��Y�W,�KYeu�BY{Y����H���/�����}2M�; ?9Pjp���Ă�tTL��\�v�!�`�(i3`�U+�PAc��N�wC�����էam�XR���b�>��;C@����sђN�1�c��N�w�Q^�MY:��Ok��@����9��;C@������Jl�y0[����	��N�Ae�#�k/�z�xEQN�By3��<�]�!����M[��ǢR�����N�By3��<�]�!����M[��ǢK�h-L���H�B���5�¬����"���������5	���]���>����C���N�T?w�����5	���]���c�A�L'Qī�*pY��am��	t���o����s����Z�n��[��{_8�Y��=�}�Vݨ�,bxqX�a���C154�EY�o\��]KOӺ�
�M�����|g�Y�'���Xw�P���w��:
1���Ƭ����
L'���Xw�P���w�S=e�d^�a��|g�Y�'���Xw�P���w����p���|g�Y�'���Xw�P���w�>0�֠��|g�Y�'���Xw�j�7���I,�D�y:#9�]�B��`6�����������s���,0=]^	�&xY�J��ev�mS��0M��y��I�+��T���jB�Fg�Y씤`��p�܂aQ�"6�l�:��h &�=pe��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcq�P ڨ�| c�]h�۟�r�@m��+�<4��ˌ�ň��h��]�F���������:C�-��5����`K?�},�F'(̺���j�e�c5���\�v�>X��ꔘ}�
�?��@�/�.��B��+ H=]A��O�T�ҹ'-�=l�)��%�� 	��k��#��5MʶE ����0*@$`��)^�T�H����d�٣��v_���Zo�����]��O�M:R	�G�L3cfi����hD�v�l�Ū�TD���)T&I2WM�vT�V��|�������c�A�L'��~�2�?�B���N�gl��ܬa(􆿳���2����.��DP֞ E2�DZ���PZ��8��"�7�r�S�ML�[�=�5x�����Y$�����+�J���q���U��@����gG�Jh��q-�Ql��u�7s�9���o>��l%i�-ݓ��E���¤�<T�<�gq}��Z鎬�������(����F�dH�/�R��(�ߜ1�D�P�E6����dE���un)�s�ި�b!��u�"��
"�,�>E���]�!����w�Հ㊟�߳�wM��2Dg�Ĳ��+�J���q���U��@����gG�g��t��ʻ�(%�7s�9���o��S8�P?_������`y����@����gG�j2��q���Ok~�7s�9���o>��l%i�-�
�CӞD��������8�S_&Z鎬������_�,�9�+�\�:�.�N��&�ˮ#��Gό���.�}�
�?���U�R�ܬ�mо�d�٣���N N�S����o}�֡��(L�^5зq8�Ј'���Xw���,D4�ɯ�U�!�`�(i3l0��F��jBo�A;h�F#"�G�����G�����!��'�(n����Z #��S���N|}	�����(S���Lp��i��F�H	5Ӡlf��`�j`������Q�DxޅR"%�ٛ�`�ί�k�6
�@���"��y ?����O�R��)t��5���p���F�!�� <&�M#���}�|f@�x�OC%��gG62WY%T��BP#�I`��;C@����b�/�J�m�x��Gr����&y�p�m~|���S�o�h<�7�ܥ��2�`8�Ȼvr��f��p�b�z'hۉ)�E�`����)��͵avF�Fď�~�26��\�eK&��s�7s�9���o��S8�)qcA����ih�b�W��{q3���y�3�!���{��~�26��\ '��O�57s�9���o��S8�)qcA�����Je}����,H/�� ��b�FP&����҅x�]�V��qP��*ӸyO�E���%�;���EWr�A����[�]�!��	Ǹ�y85�90A!*9�5�����Ƀ�.��|ȃ��p9�"3�ˈ��1���J�M�����y��j��k�G�ı�!��"� +}���k$ mxgQ�3\M�aW���^��^ٵL�wy<ڃAH�RtV�^��vf�<�R�{_8�Y��.��ib��}Dq�f�1���~��$o���l|�*"k����br�#������0�	1G����sC���X���y��lD%~V�qM�)FŒ�J7
i�c�r��5ߧE4���g��A�uۥ�w�BAGeG�3אY�{'%s2�ew�rcF���;f���Ն gWVbT+�q�7B�[��(��� �����W4%��!��z�."�)��5�-�B�7q�|����ʷ5��.�U�
{�~jTK��>�scX{�X!,G�&ց�*���,픿�n���}���S.�3��)P<�ܓ�Y!�`�(i3pı��0��ho�����Z��3��w��\�W��?D�8��ݓ�W���o�0�\G�4�0 L?ஹ�%���M�Z哚��ݚ�Н�(*�O�q����j��[}�N�`2���K��K�u�>>!�`�(i3�[<��؅�&~e�e��E{��h�^��x�`g���|e"ʁ���MյvϬ��	Ղ�I8�y\��S��z�-G����|!�`�(i3U /숇��"�ܸ-�;S5b	��T�.�N�h�9���6��4�2�|�A��U젩`#FW8�	���:��$�8���}Dq�f�G�&ց�*�=��L�j�\n���}���S.�3��LX�N,S0!�`�(i3pı��0������X,�Z��3��w��\�W݇�g����ݓ�W����bh�UUd4�0 L?ஹ�%��H~x�l��V�ݚ�Н�(*�O�q
��O���[}�N�`2���K��O_�	�b(U!�`�(i3X+�{`����&~e�e��E{��h6]F�#S-���|e"ʁ���Mյ����J4��	Ղ�I8�y\��S��z��,fף��!�`�(i3U /숇́�y�62@-�;S5b	��T�.Ϧ�R�E����6����r~�4`��U젩`#FW8�	�����W��bP��}Dq�f�G�&ց�*��a�	K��n���}���S.�3��d~k�7ZyM!�`�(i3��O���b�z'hۉ)�Z��3��w��\�WݯS���HN��R���
�Ŏ��HN��R��Gu�"�0�ʥ�nr] ����h����zNc5��;�P�t�5��f���,hʢ!�5��=l�U�-V��_?i8qE��6I&���#�B�k�'y�/$�ߺ��]��T)��>֯���,�*�F��cny��&�;a"��0�혅vº��żפ	�?9Pjp��17e��:r����ZqJ?�d���&��ꢤ�Og1����?���zf�l�=U�0��IuAv/fu����1��� �U��֜��3,0=]^	�&���忑������Ho��'�\�n���D)9W ����,�ǰ	M,��rER��?إ�c��Nz�ً��:+ᕺ!�o��φ��<�6�$>ʹ�*�Ĺk\������`�5Ԍ������@�:t''W��Q�jI��Ͼ��\]�Y���v�岦�%I^:��%9&���;���EWrqi}�Еi"�,�>E���2,��T���$�Qu���(��h�)�W�=�k�i3<�f�D.`�Z���N}�m��{��{&<c�yQ���4�5������-"{b���~�26��\x`]N�~!�`�(i37�ܥ��2�'k��� �&�C�|检+�9�jɲ�1��� ����P�7� 1�ж� �4���܂��+x�r�u�#��nt5޵3{�aP�E����F[s�9�-n���~�2�?�B�����lC��U�T�\ ��yO�E���%�;���EWr~��*i"�,�>E��ʆ�In��t�8&���I���8|F�KD�Vr[/}>5��0�B� �b���H����o�γ�ha��o���H�RtV�^7O�D��w��N�Cٺ��#o�]�ʄ��.�L��w)��
=I/��\]� h�ҩεSENan&���ߊ�ֲ���ܜ?n昼�2#:�^�V]��}>�C�;�����:=����l������6z:�B����]��V����l���.�et�rZ�?ђ��P^(�՘�}���������J�\���=��}���)��U�UH�RtV�^!�`�(i3z���r#� ?����6	�T��u~��t����>PQ%cp��g�H���~��!�`�(i3���F1������$��\R�j°��ݚ�Н��Ra])n#����0�������ߺ��8�ۦ�P�X��P�������pC-��h�:�	4}�sv�{��qWU���>
A��%��WG���;� h�ҩ�!�`�(i3k�s�X�C�GM��4�ūd���8tO�M:R	�@tqx���!�`�(i3`
 ֢��؜J��v�S1��6�uE9�+��!�`�(i3����١�$�ݛ5�CNi~�N,7tL���4X%��C_=A�H�RtV�^!�`�(i3
Cj�R[z�(�� '�i�*ڃ݂S�����3�t�.K��ߎ�x��y��v�9��!�`�(i31}�ั):9��tf��!
Cj�R[z�!�`_q�!�`�(i3�̢k����J�\���=��}���*rcxm�N�e�{�W!�`�(i3h큈���g�W����w:�눔�C.�u�X��I�ՠ��t����>PQ%cp��g�H���~��!�`�(i3���F1������$��P"G�wk��=MNԅ,+��}Dq�f����%>�rGO�D mWN!�`�(i3��֖+�){?a� ~>>ը܅%GbNÌ�Y,�u��r��!�`�(i31٥xu5=�Р��U�1Q�\��^����!�`�(i3�	��x��ݚ�Н�����l�鉌(*$ΐI�q����!�`�(i3c���P�vћv\���7��{����S����9�@��!�`�(i3`
 ֢��؜J��vv��v�K���x����VY�l��NI��ݚ�Н�
�:qEp�;�P�t�5!�`�(i3$f��_Ub�F�S�1 �fĉ>99��R�Q���~��p�������l���7�����Vq�|`kK��I� zSd��;��-����!�`�(i31٥xu5=�Р��U�1Q�\��^����!�`�(i3��Ě�����}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���ء�I��߸��S�Ȍ'�� ��@O�wR��_��3cה����:
1�������t�T�s��"��;���EWr�P�SYG�_�����7k��/j�Ch��㉊���;���EWr�c�Em��W0i��^��{��e�ֱ�q���GH�r@�Wٶ���3p��Op�ե[�u�,�s����+�^n=\f�5>��kV��ܜ֯���,K�~��B�0M�Ŷ�Eʨ�`N/������&G���lS���|�+^/�����������p"3?K�[<�6�Q=�U�E�0��0?�R��e�E��4�T}�Y�PG�(��"��&H] ID��RN�1��-��	����#����qk6�<�Td��M�/�}���[�L{���k0'��Uo�� 
r�16��,��/�}���ļ_)a�0��-��������&���:
1���Ƴ��d�L����|e"��jVѭ@����&���:
1�����#QSU:�����|e"�錐�� ��M��,�4����*~�ݚ�Н���=�g[V��M*?�},�F'(̺���=c��� ��Q?M8�f2!�`�(i3����*c�:�3���nu4Bޗ��;�fޟA'�
�:qEpCt�w#��@�ݚ�Н����F��O��;b�-�2��;�P�t�5�{�6�C������n/��dc�@c�����h!��"� +}���k$ 	�!Wn"��/�}���ļ_)a�0��-����m�����GI����ht��ܜ�[�״$(�>g�������'{w#/ B����&���:
1���Ƴ��d�L����|e"u)^��r�Sŗ�}m<�{�6�C������n/��dc�@c�����h�E�i�m}6O�D mWN��ܐ�}�~(����[��l�,*���E�D��Y��<���y��,���o��_�Rv�䩲$����E)e|A��`���φ��<�6�B���ؐ1nk��|n�xjzӝ���w3��׍�&�U��f�P#+_]ݱ�p-����`�(]�`��my$�N��o�/���;�̢k���F�KD�Vr[/}>5��0�B� �b���H����o�γ�ha��o���H�RtV�^}I�6����!�qgy�`��vN	���QC�íN=]b~*��s�)��7��Y( z�P��1tSjv��B�'��a��¤�<T5џ�<)@ Nf��#zP!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN��Ě���aT��3G�IX0F�M� ���Ī#e��K�� ���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}ڭ�X�Ә������Me� F��pcew��y%>��˳�Ş��"m����f���Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�bƑ��'lv� �0#φ��<�6����pIy��$�Qu�F��&�o�WW;��'n�^0o**�ХM
�nGZ��JP��(�ߜ1����˟y{y����i�q,?5qj�����)�E�SI�k��Xmt�=���3��a���!@�f")u��r���5>������y�!��_��0J�M�����0�9&،��F�z�8#Ҟ�#�>�L��n��p��b�Bϱ��>1J���ƈ5$YaV�Ra])n#���r������N�T?w��OZ|��������Y�I����Ě����DU�Y�K��
��
jY�o�v-7�I�q����!�`�(i3V��N�xֳ;F+��]�����4��.}�՜�D��s�hX�ɣC�7�/�)hϬ#�gnA"�߿�wW���Z<��A!&�2����M���CO|e��߬�x#=���c���9���G��+tt��H�����}�tץ���q�H��{���U���C���C�7�/�)hϬ#�gnA"�����ӹ�Z<��A!&�2����M���CO|e��߬�x#=���c���9���G��+tt��]�3��=9tץ���q�H��{���U���C���C�7�/�)h���Я Y;�Uʮ�V(Y6� f$C�{���s�y��j��k$>"A��⸱n�����?��#b�.]����q놕
�w�m����fh����p���3�eO��W���[��l_�0\� ��+U���Rj:;bK���ţ��N����������y�m|^�XlF��%�K�7��C����)�����iZ��c�ڭbK���š�e���L����$73�E�eNzL�lS��V0���w&�.��;�P�t�5HN��R���ء�I��߸��S�Ȍj�����)�n��;,��6<����G>6�x�Z2r�D���0��XJYOݸ��-�eH�4)��U��)���Y;e�iK-pm!9�>��n4s1�U��B��-���N\�͝�!����7�癆cgR������������ h�ҩΡ�ΐ���-a0a3�8���[{/;k+Q�h'�Ȝx�5W ��̫(� h�ҩ�:
��x�{�\��N�Ś�-����;�jmT�#P���1; ź��p&�{�A.�<���H1tSjv�
�:qEp͘D5��'�^�����ݚ�Н����F��O��ݚ�Н��K�,ǆ�`�íN=]b~*��s�/$�ߺ��]���޵.�ۃVa�ir=5.B�����'����u��r��tl�:�K���(L�^5%��v��!�`�(i3�5ߧE4��
�:qEp�;�P�t�5$f��_Ub���uQL+��φ��<�6���ΐ��S����N��/Z�o���vP8ԍТ���hM(�s�;{����B��ҧ4�@	�u�a�ݚ�Н�!�`�(i3P�j����9��"<\�}
T�W����9�kҦ�!�`�(i3!�`�(i3!�`�(i3��jVѭ@!�`�(i3�2 /��u���3om���U�R^p���P#�w�����U�R�ܬ�mоf1�.��N����k$ !�`�(i3��>)����E"�N>I�AS��0+K���t�T��?E-h���U���e��_	�Ƽ��S�J\70C.�>��V�m^݆��xjzӝ���w3��׍�&�U��f�����C؆�1�u:�3u��b+}y[�k��^�1��dc�@c�����h��-�����s�Yls�<Ԍj��_�mS8<�n�ݚ�Н��K�,ǆ�`�íN=]b~*��s�/$�ߺ��]���޵.�ۃVa�ir=5.B�����'����u��r�����C؆�1�u:�3u�"��ӌ�r���%>�rGO�D mWN;�jmT�#�0M�Ŷ�Eʨ�`N/��R��3���:
1���Ư����z���!*��*8b�3��_�mS8<�n�ݚ�Н�� �@[�鋽C�H�CW���|e"$f��_Ub�F�S�1 ����F��O�}�	76�&�� Ӗ�t$�)�vxj�y��j}������v[2�quA0�e]'\gWg��	�Z�kfcj��r���iI9�o«IX0F�M�p�	�\���F�`y������T�8k��.ͥ�H�RtV�^�N�*��	@n��뾦��߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#��"����G��Hb� h�ҩ� ���Aؠe
�M����d��-��!g��J�s��z�
1���;#o�]�ʄ�k�q@g����Z<��A!��-����!�`�(i3�N�*��	@n��뾦�!�`�(i3�5ߧE4��!�`�(i3[�5���78�íN=]b~*��s�/$�ߺ��]���޵.�ۃVa�ir=5.B����<���H1tSjv�%?gV��Ux	���G)P<�ܓ�Y
�:qEp�;�P�t�5fĉ>99��A0ok�����F��O�\E�W��4bƗy�"c̜�&�f��ǩh\K�5~�0��=�e
B%~��6�^�z�@��E��?J��W��x��[=�zɣ��S`&c�'N�jX���˫φ��<�6�@a� ����C�'�ąd�G}%����3f�Ȝ��Y��!%9�G�C\���F�`y������T�8k��.ͥ�H�RtV�^s�Uo���ַ�����ƍ2���l�����g�Z��3��a���!@�f")u��r��$XR�QܛOcOZail������&G����l�� ��5%q���f�e�x��w�����q� Pʬ�J������nT�j���c��1tSjv�V�Ո���߿�wW������4Yz����|e"$f��_Ub�F�S�1 �6�>�@�	I\��Y� z�P��1tSjv�V�Ո���߿�wW��C�H�CW���|e"$f��_Ub�F�S�1 ����F��O�}�	76�&�� Ӗ�t$�)�vx�m`����Z��b���Q>�<��#b�8��B�5�¹�*��a"N����#�T������oj������ZN����6�o8:4�I���c�90Mj�dL��~�26��\;��B�lXm��G��*IÙ=�HV%~YqsوiI9�o«IX0F�Ms�Uo����=Djw�9�xjzӝ���w3��׍�&�U��f�Dw\����ō܈��VW �+��!��"� +}0�ʂ�j�Ï��	�l�lM�3 H�RtV�^L�J)���� \L�1tSjv�;�jmT�#V�I>1͊���3-��g�MSG~1tSjv�!�`�(i3�����i�X�-e/p���C.�u�X��I�ՠ������&w`C����"�:5A��p�	��x��ݚ�Н�Z��JP���K���&�9�ڟ,AX3�T�#_�B�ݚ�Н�HN��R��bP�63Z�t����l�� ��5%q���f�e�x��w����֯���,mk��L��wd����s3��0��"(]��� z�P���T�ݡp��b�W�
�~�m5�)C�]�Լ�c���J����ݲt˻=�}���yb���XUIl]��u��r��Dw\����ō܈��V��*�f;��}Dq�f���Ě�����}Dq�f�Ql4�ul{�]&"(�'����u��r��Dw\����ō܈��VW �+��}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���ء�I��߸��S�Ȍ-�+���5FY��:�m�91�ŴbK����֭�wu3���l��
��Mx_��9���I�)+��������� �"ƾ��gx�׈�xIY��8>h�|�Ȝ��quA0�e]'\gWg��	�Z�kfcM��fZ� ��b�FP&��N�T?w�W�E<HӍ��XP���ʥ�n2`q:Fa�7���⾰��bK���Ŷ�����\���F�`y������T�8k��.ͥ�H�RtV�^�Uʮ�V(Y�t���1�g)P<�ܓ�Y�̢k���F�KD�Vr[/}>5��0�B� �b���H����o�γ�ha��o���H�RtV�^(܆�NGV��}��6�8�-Zy?X���a��ݚ�Н��GI�\�0�c��v�'�i�*ڶ�UKs,��#��I2�8� S������v�9�ʒ	��x��ݚ�Н��GI�\�0�c��v�B^`ٌ���M���
�:qEp�;�P�t�5����l���Оt=�[&��0�|섃Va�ir[��l�,t���H[W?x��w����]�Լ�c�#o�]�ʄ�}�V����N�T?w2Rԟ��n1tSjv�X�o|3bK�����`���UK�"��ӌ�r���%>�rGO�D mWN;�jmT�#��U�R^p���P#G��Hb� h�ҩ���೹�C�A�IS��[;\v�a��ƍ2���l�HN��R��bP�63Z�t��Ě����E�i�m}6O�D mWN��ܐ�}����L�yE�:�.�N��������m>�G���'���V&H� FMsO�~�fB��t|ql�osZp�W���
�$������%H��|���2,bK��������H���U��)���Y;e�iK-pm!9�>ֱ�q�����ѧv;�?�@,��VJHn��z��r9�3d�G}%����3f���L�yE�:�.�N�������a��r$ɓǉ�.y�U=������&G��೹�C�A�IS��ַ�����ƍ2���l�����g�Z��3��a���!@�f")u��r��$XR�QܛOcOZail������&G����l�鑴HH��"�̙	,N��>�s�,�H��-����!�`�(i3}���yb���}�@���_rS�b�8Z�AԢ�a\�2}$#h6������t�_��ݚ�Н���jVѭ@!�`�(i3}���yb��-H��.�����o�����[��l_HN��R��bP�63Z�t��#�a�Ą�ԬQ����5��t�	���QC�꠼*d�m�d��-��!g��J�s��,ܓh�,�;�W�m�-�m����dBu��r��a�}�$�᢯��0���O|������NM���fĉ>99��A0ok���H�����Uʮ�V(YhV|_��a��o���H�RtV�^w-)Sz�MB~�S;���C�H�CW���|e"$f��_Ub�F�S�1 ����F��O�}�	76�&�� Ӗ�t$�)�vxկz|h,�`_�o�@^¬P�ChYB!c�3Nφ��<�6�@a� ����C�'�ą�2N��n��bcb�q�\�K���&���\�v��_�R�G���+�^n=\f�5>�yk���]{�7�癆cgR������������ h�ҩ��j<��?��;c���k+Q�h'�Ȝx�5W ��̫(� h�ҩ�:
��x�{�\��N�Ś�-����;�jmT�#V�I>1͊���3-��g�MSG~1tSjv��0�9&،��F�z�8#Ҟ�#�>�L��n��p��b�Bϱ��>1J���ƈ5$YaV!�`�(i31���~�0�9&،��F�z�8#iY�g��Ѻ�&\VI`,"#S�K�.�$f��_Ub�F�S�1 � ���Aؠe
�M����d��-��!g��J�s��z�
1���;G��Hb� h�ҩ��H����ӔРq
V2?�@,��V�=aS�H��ݚ�Н�U�z���K� |�>�!�`�(i3��jVѭ@!�`�(i3u�st�⫴�IV�*F/��}Dq�f�HN��R��bP�63Z�t;�jmT�#��ΐ��UG�*"�!*��*8M*QfY�"Z�';��#j�ݚ�Н�U�z���K� |�>�!�`�(i3���F��O��ݚ�Н����F��O��ݚ�Н��k��M��5ߧE4��HN��R���ء�I��߸��S�Ȍ��̓-��w�T� �f&���#��uގF1he��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc!N�'�y�G