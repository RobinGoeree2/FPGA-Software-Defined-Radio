��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���G�H�ƻ	�"�iQ�����3�7Q��㼫F|�ݽ0��@h ���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�����|"3�����U���T��ײ2��>���^k�/7�?1�(�c��ߘ�]�~"ɟ�S��P�jh�I�?g�f&:��r-,�Ny5�7\F���r��C>C�݂�N$��/���	�0���'v6�o����"���Vv��x�۔7�D��:�b�#�Bn�K�͎��uP!ߌ��˼�{�&��,h;2���۟�
$�e
�9��Ax!P����Oy���9����^G��5 ������2Ee�Y�R2
�I.��	���
���s}��=M���c���X6(!2��탯;\߰`���n�T�ƫ���7 � ��"�!Z�*_#a�|�82�WF�bK�'F��������)���UeB�G�g�vvS�}$�SK�m2I=������$�
�K�Y���p��}�ֻyޟe`�m*]���G_��Z�x>x���N�/ ����l�Bk�FB}��O5rQ^5�y�0+;4ڝ���&	q} �<� C��\�'uOe�[byPN�pj���Ʀ�?�¿�b��T�Q5�P1aq�q*�{������gLE�zϼ=�Db妘=��"D�cHF��eUٻo���mi��*	�ť�.^�i��' 1wH�x�xs��3�<A��z����
a�������~�+��,/,����W >g1�]l�&Y��F}갨y�����# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��`y��f2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�}�Z���ik2)�
}wʭU&H�1��8�h7H�u�ÍeRuw�C?3d,f$�7Q0�"<�F�ٴB�I�SbW�'f�ٵ�lf)@̲#;���(�s�-���f�i\􁗊�n��\v;V[���b�/Qk�� h���Bzb;ym��+a��ʁކ�+��T��C�NJ���1�:�Ω�*���g S��/P�pݒW*g;X��'p�@�I�?g�f&:��r-,"�却G�Ct�z&��ÃlO ܅d:��+���������i�����X=n/a�τ,HKObM�^�T��a⨯�T�w�����.��֞�������i�����X=n/a�τ,ʨ�lC!�!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�{���exL(�M#"�?L���u�p$���"��SM0.�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�XW�������P��Y��5�d���I�'z�Y�f��4V�H�%��F��F\L/���?T�=�4e=��-�ĕ|G���!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3.N�DMY����U��t��ܣ^\t�*�00/ 	CH�.�!�`�(i3!�`�(i3!�`�(i3!�`�(i3���y��lDAͨY��ژ7^2$S�6���f�����C�!�`�(i3!�`�(i3!�`�(i3!�`�(i3���y��lDjg���֛�:̚�Fu7V�Y�\Jm��MV� c�!�`�(i3!�`�(i3!�`�(i3!�`�(i3��}>Ό@^�����4];ˍH����D��ܒ}�X֗�P3z}�&�!�`�(i3!�`�(i3!�`�(i3!�`�(i3����j��L*.>�+k(a��H�;Q��G�S>$XW��WA{I�Z�T�����N��}Dq�f�!�`�(i3!�`�(i3!�`�(i3!�`�(i3R���Xc���a��_�`��H�I��E��4�T}�Ĉ������=���f.K!�`�(i3!�`�(i3!�`�(i3!�`�(i3Ta�F�O���^�#��\�'k(a��H�;��\_9ͫ�}	�WA{I�Z�T�����N5y���=.���'{���*��O�t;e���`���ҕH{6��!�W��!�`�(i3!�`�(i3!�`�(i3!�`�(i3Y�4Eb�������犡�&Y��V�5.Pf����#�u�'�'�7��r�=!�`�(i3c��Et��q���U�ЂDa��(o��0��7�E����F��j��\w��0]%��C���B��+ H�����5	���]���[�(>5:��f�C��Ʈ+ˀavM�)��� �@��&}!�`�(i3N�By3��<�]�!��	Ǹ�y85��3}�@�7"j���b7|#9���{k�h�+_���&#ݟ�"B��$I��w��,c�A�L'�����CyW�f�t<|������N�?�_uM��y��I�+��T�����D3���t�  ",��%���E�EYZ/�矘��-n��I�?g�f&:��r-,"�却G�{�.���qcW�(u�" Oag�֠$b#^M�Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�t�|�Q�(����ޏ����\�'�o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��c����^b�%@�c�3稨�;�}���-�Tu+J�����iА����H�Kc���- ��5�}�]����8�z�G���S��ȯ�By�`�2*Q=F�k�mD#V���)���6��,ڒ�p��e"5�O�%E#P �s9r6�$;��l�6�Ύ)�VpPOxtX+�YrM�e<�Z���L`'���Xw�j�7���5�%]���a(􆿳����^��b!��u�B��C8�4a��!����  ���d�G}%��Ď��J�;փ�����ɇV�"S�|�\9S�l���r���d�u�׽%��]����7|)�` ��%J%����=� ò'�����7y���;6٫�e��nb�� :�Kn��u������^"�p��ν(C�|�R�n*R'��#t��s�bМ���yU]�����t�T��?E-h��$^(?��"��h��w���`���φ��<�6�b�� �I2�?W��z\���F�`yx�>�+X�[�G���K!�`�(i3<�6�Q=��S<����K��!L��3w #�T�Z��&�2������E/��F����R gWVbT+^���1i�7�N��i���:=M`�K)��v�^J�&t��b_X�XV�b�z'hۉ)��d�7�qĉ��%>�rG�E`���՝� s�#0�ʂ�j�Ï��	�l�lM�3 zM#��m�.�
9� ���(ٗ.;��
�6�j�<�6�Q=2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��َm(5�X �^�(�R��W0�	�:]IKp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��OC�0����l����� �'����u��r�����voȠM���¡y p)2ߓ&?4A�5I��!�`�(i3C���6YU�ǔ���<�
�d���ƒ����Ș&����Yk�����voȠM���¡^aE,K9�M���¡�ǳ��&�!�`�(i3fF�5.]����}Dq�f���Ě���ž_�F����F��O�}�	76�&�φ��<�6�b�� �I
SF�=�g�{k�h�+�_�E=x��M���¡ȯ�By�`�!Ʃ�T������,�ǰ;փ�����ɇV�"�,\�B��?2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ�e 4G�1�����{�a|����$��$��m4�ڲ�{���4�Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h$�ҞC���aD��3MA!�`�(i3!�`�(i3���Y\_�rM�e<����)����B����d�+�āK��2WI��o���-�� ]~T2��4��)�Bi�v�Vȡ�&Y��V��ۋ�8�u+h���}둮�Z�)��;_�O+��B;��|B��� OD���S��ϗ¾IŌLNk�#��ϸ��#|ShI�ˋ��X:��+�<6��$)K!�`�(i3�E����F�׈PzO�e�n�^�(��.��dLG���6!�`�(i3����X=��}DD����}Dq�f��~ fbܢ�{㯲��!�`�(i3;/�"���_�����ݚ�Н�Q��=� �9��X��ŀ�!�`�(i3�:ET֤vKN��B�)Y!�`�(i3?�!�`�(i3!�`�(i3��TG���P ��*��Q���ǖ�!p����nZ8�����
P=ܽl.��n��s!�`�(i3�E����F7G#+�Ǘ0z�cUL�2�c�L��lC��U�T�\ ���:5A��p4���v�d�!�`�(i3!�`�(i3N�By3��<�]�!����M[��Ǣ,�ttT��Q�#<4^�!�`�(i3�����5	���]���>����C�=�M����FfL!�`�(i3�����E��@IE�U����S8�gY��U�v���W��_�ړ8���/���}Dq�f���zsqG�zM#��m�!�`�(i3v�ј�"��Z鎬�������(���	t�����"j���b7xY�J�����ǖ�!}�	76�&�e�0
A���W���b�0�� VU+I�j.$�)�PM�^-q;6aJVlO/�ݚ�Н�b��
ߎ� n2ϒ�ȡ�&Y��V�
�V_nu�$�F5k0B�����l�����\��w��;���_���	ލL/���?T�%��^[�r����'��,#�@�΁�a�n���l�|���jWɆ&6�\]1]�?���(��.��/��lӹ��zigzA=v)����X=��}DD����}Dq�f��$�V��bst�N���!�`�(i3;/�"�����h��!�`�(i3��5@~Ju*k`Ë��!�`�(i3��TG���P��7U��s#2\z��}�� �с�'(�U�c"�,�>E���	h��IB��`���o�?X}Ax���x��~iM5/�S3 <�E����F�׈PzO�e�n�^�FR�6�!��&t�ND��������X=��}DD����}Dq�f�%Y3(�6��B�r��!�`�(i3;/�"��ZdN�ɁRN�]�5'��}Dq�f� �	{��/��@����^�v�!�`�(i3"�,�>E����-��%Mό���.�!�`�(i3եa�����!�`�(i3!�`�(i3c��Et��q���U��ݚ�Н��AO !�`�(i3!�`�(i3�����
L'���Xwd�n]NْJם����"X��[��Q[R�7`
 ֢��-�¾L��!�`�(i3�E����F��j��\w��0]�wӨj]h�u.$���!�`�(i3"�,�>E����-��%M�rs�i�نW0��;�¬pX��g��U-�e oȍ�~�/���i� �B0��O2��p-!]�P9d^\'@�6���{6y
N֜�s�b9������|L�K���3P�|�2*Q=F�k�mD#V}�D8ҬϦ^c!�6��[��l_�5����`K�o�f�ԜǄ		c�S=�4e=��-tE��gV��tR�/p�ΰ����4V�H�%W������\o�LCd�,��yH��!�`�(i3���+�J��Y�{'%s�Ǹ2���;�¬pX��g��U-�e6R��h��˽0?�.���J�LQ��wb!��u�C�m�n!�`�(i3�n`5�fK��0z�cUL��Jv(K�V��W��_�ړ8���/�I;��3�>{j&:����SM0.�ݓ��E�fZ�z9�Y_䈵v�q��T�ٮ|�,
�����j������Q�z8!Ǩg��U-�e�,���6+��n~�x��&��+������ꀍ7s�9���o�jƓ�[���+�^��BY�B����葏���͸|t��R�
��>�.�C`S�r5�ۢ�2*Q=F�k�mD#Vֶ�������F�cZ��K��2WIK�d�rM�e<�:v���Z���d���!iO.C�+��uK[F���,!��_��Tq�'?���r����l���r��|-I@��v?&�2�X�|������r����o����D6�~�ݵ|��*뇮� л����U�p��X
�S�9�\%��V*_�ِ�b0Q���$VǽO�~���c�.��.�rý�5s���Z��g St�T�φ��<�6�@a� ���N���Q'݀�=��`���φ��<�6�&@?Y�#y�vNd�)i���"sS<�0�zG����ZAL�:!�`�(i3�d���a؅q$��.��m�f.���G�?v��� �+��R��!�`�(i3¤Gh2�&x����E2b�z'hۉ)��d�7�q�՝� s�#0�ʂ�j�Ï��	�l�lM�3 S��(8n���ž�Ć�T���7X���c�}��H����o�γ�ha��o���H�RtV�^.�`��ai��ΊqE�?4A�5I��!�`�(i3��Ě�����}Dq�f���Ě�����}Dq�f���ܐ�}�۪�G�;��O�I��)���W�w��fD���ӽ~���Y�b��K��*�:�b��t��0�$�Dd�V�E	��J�6�D�jOs)l໶�,!�`�(i3!�`�(i3!�`�(i3{\���!����Y �6�$�<���U\���� ��\_9ͫS�# [�T6�`g��Ȇ�k��vy�eč�0P�{��d���!i�Ѳ��a�\�2��3-N6����L~�4�����}��`��GedTly�)��)�`�(�@3l|�gV��r��B�"}��o�u�/�tL"[$��SE���� .[^Cf|�9���������=R�b������'��8���f}o�Õu�RV��,�X��4tΘ�2�9����럍�IJ�� ޘ_�92j�`$|˂�I����,8D���,=
��P��bG�d8;¯C>��Ӛ|s�g*n{�Cy;"-���n�|�_��Tq�'?���r������o�	�=��Y�$���E�i�m}66j�"Hs��^fp�/~ �GG.�L�7&o����@�\�FUX�u��ȋ�=�^�Na�gN�3c!�`�(i3!�`�(i3!�`�(i3��mqf��x����y�mZH֫&]9�(b���J��:�������+�^��BY�BAsr�7���X�u��ȋ�=�^�Ny���0ܔ������*[wL>r~�/����ȤOa�u��KZKQ��G�S>t�:Nf�󑾲YT&9.��o�2L;���x9;*A���.~0�
n���68;�
4p݅.�g3Z�)V��B�1W���.1	Rv�_�-6�v'���@P��k����Q��w�п?G����C!�`�(i3!�`�(i3!�`�(i3�����,��gCu(o?C*
��10�xJ��:�������+�^��BY�BAsr�7���X�u��ȋ�=�^�Ny���0ܔ������*[wL>r~�/����ȤO�����l)�F��A3-���X4��׹!X�%c�3p�dr������=��]�w9"x{��R�w}�	76�&�;��|B^%^0��j�f����3a�.`Z�WN)� ��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�ƹ9��Pd���	��B�Mt.K8�����葏_����B�!V�����τ~����p���`�D���)�+��u)����w&lO	"����-{n�͆�J��!fWUVƌ��]�u�|ʓ����k9?�\�N!V�������F$0y�ׂ�G�3>q��X� 2�2��Ȅ&N�b�����v����5E�Ra+�u\ޫ�r�$^���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc9g�O��B~&�ȫqO8uDb�G�r�y
N֜�s�Y��"��5�O�%E#Pd�G}%��Ď��J�'�J:��XDf5a�҉]��H��>/Bj�Ւ{K4P7�#�'lo<��G�s2F\�M�M���bF��ϸ��#|S������3[�u8�(��.����ֈS�&I=�S��M�����H���x!�`�(i3�$�V��bst�N���@��?\K��i�ڿ�ቬF�Ԥ�5=9��n�7�Y��ݫ�QSV��� N"�0�i.�9�
P=ܽl 6�+��(��S�t�bS��L��,0���\N�A�~�Y���(�\w��B���t$Q���31�P�V�!�`�(i3�k�O�>��+qѭ�+g[�!�`�(i3��-pө[��&8�,�r��]����f�?ǉ�=,�ttT��Q�#<4^�Tl�������l6�=�M����e��F8�D���K^�)ӭ�r�#U�!�`�(i3=�p�N�L�!�`�(i3C���VK	�)�^�\?�)�O�8�W ��A��X;p`���y�v;�RN�]�5'�E�i�m}66j�"HsS�~�L.��dsBj����?��b������?9Db�G�r�y
N֜�s�L�-f���5�O�%E#Pd�G}%��Ď��J�Tm�v��G��G-"ұ�����*y}e�^X��4Yuc*�uM��%�p@!�`�(i3�@U��0�To���.͖�:�U���6j�"Hs`�0�$!�9l��b�[�N5(+Wp�ΰ��QB,�<�>_��X'U���P��\_9ͫS�# [�T6;��|B'O�d��FiI9�o�?�d���&�8���SY�N��j����g�o�3����"��є��&Y��V���J�=@�%��j����Y�4Eb���I!����)��Uza?Yƨ@0�$��ѯ���Z¿i!��j9'K}+�a�����'�u�ȓM�Me��'�ZX^�O�<KҽX:H�RtV�^�Ǩ@�z�.��"�]'\gWg��	�Z�kfc��2���8O.C�U��B��-� �ѕC?"���xя��!�`�(i3�'ž1�|�'����z.��W��!�`�(i3NL�Sfo�r��n�"��Wr���,(��9�e���}��2��}��D�o�&x����E2b�z'hۉ)��d�7�q�՝� s�#0�ʂ�j�Ï��	�l�lM�3 S��(8n���ž�Ć�T���7X���c�}��H����o�γ�ha��o���H�RtV�^;�jmT�#⼲Y��pJ�V�G��Hb� h�ҩ�!�`�(i3p�n��E�g�������(ӈ���m�r����!�`�(i3��jVѭ@!�`�(i3q�\E��0d<��2:�OpkҰ$!�`�(i3HN��R��bP�63Z�t���%>�rGO�D mWN���%>�rGO�D mWNHN��R���IX0F�M�Ǩ@�Ws��h�G����,�ǰ� Ϳ�&�v_��Tq�'?�Y^y�*ܦ�i��>��Қ�"<T\ �r,G�W�"�Ů7�6��,�,�W�8"M�5�O�%E#Pd�G}%��Ď��J� ���骊
|�g.��g��Gt�{#	�x�7M	�\�4���u�vp�$9��K�Q&��+���Qw�c4~Nrާ�����ݚ�Н�!�`�(i3�~�7p����nt=:�$r�t�}iV��	��y4��$�[��{8_��h"�+�r���)`s﫱Och�����ƛ����0�^�!�`�(i3!�`�(i3!�`�(i3�����,��2*Q=F���q/���<]9�(b���J��:�������+�^��BY�BAsr�7���X�u��ȋ�=�^�N�˧�h��.���L2��500q~I��aFN�Ң�,�\�,[����<o�Ĝ
�Y�M-���YT&9.��o�2L;���x9;*A���.~0�
n���68;�
4p݅.�g3Z�)V��B�1W���.1	Rv�_�-��*rqg�o�3����"��є���;�����]����`t1�-OY���B���)����7c�l����[ߦ^Cg��)i�xx�j�GWw�;_��]}� GK��� ���*5�$�Ƣ�/����3Vq�)����k��d���J�W�o��-���HU�����_� M/������Dݘ�� ��z����wWi:rö1M(7������C#/<���q���U�p��X
�S�9���:Y*��l�+�7#��.`L+�&�H
�D�x[u�r�S@�=�{��5�pJ�V��U��)���Y;e�iKI/B޾PԐ#��go`iI9�o«IX0F�M&�H
�D�x[u�r�S�H����Qw�c4~Nr_�mS8<�n!�`�(i3���y��lD�	Sz��
�GBQQY����#H�Yg�yi��v��BPlLO+@�=�{��5%�iq��e���b�'�^�����ݚ�Н�����湡N�Ւ>��4��yT�M30dN�<@Iv��nt=:��:5A��p*qA����6\�4�@�� �-jېI�q�������?B��#Ɵe�*|�÷�Wе !�`�(i3L�J)���� \L�1tSjv�����l��}G[���S_r������{2f�V�i��Ք1tSjv�!�`�(i3����湡N�Ւ>��4��O�#��q#��3F����Kq��R�=����M�!�`�(i3⼲Y��pJ�VҎD9��ɰ���|e"�Ra])n#���r����g����Vq���|����Lt�2�t%��v��!�`�(i3��Ě�����}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���IX0F�Mմ���4��E��$w�R���y_Nr`e���7!ךv���{Q$M�`V�����H���,>$��:?���