��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���G�H�ƻ	�"�iQ�����3�7Q��㼫F|�ݽ0��@h ���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�-Q3�YN
x��]Qu ������[���a�8%`��4�s�6�XAoeuxLZ�#8������^F��W��`��9�����u�A��c��]��;�I�����)O��Ξ4�"�\�� ���K�O�{��
2�D�� ���Jc\֣�I��B���t��|U|�/֚m� �+d��.8%D.��n�P��<2�q�U��k�8u[\E���@N1�w�0XL����[fe�Hs��9lSUQ�S��)���2Ee�Y�R2
�I.��	���
����k�������0�?�}4��ѕ�������U��=>bMab�	;4��G����a�����(�I�?g�f�P�����Q� ���6��H4�
� �AH�*��.�T�{ ��ʥX|2�
�ƴSkC	c6���i�P�GyϪ+2��?� �٠F���JlwLX�j�{~ �[D����RL�a)3���ʉ���I�_�]i�Ϗy_�Q��eD�7C��H�و�@����t����H�.�G|��k۴������\�4�si�W���jh�6g��1���5��a�@�o@���q�&��3B�Hj7�;i���D|�"G��k�8���҆�|n����5��K�O����FT��sQ6��j�'E���x��,"G�g$	~�|O���4du��w)�S�5� �7��Mv�9*���f��^(��f�)y�8�:r&@��=��$얃�rb2 �Q[1I�����w'�\�Q�3M���e�t��yn�	� �x�m��n~�q({L�51��;����'��%Ճ�86���H�aF��6��I���j�r�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�E�s��bc�Ѽ?��Q2�=W�֯�^��N�&��^˻f��	g�y���}�ZC��aNvA�;��>Oʉ��tw:g+��T��d^��_|��3g�ݜ��s8[Z�`
5��*�z�������D���J7"z��cX궘�[�nh�/;KYˆz}()pxt4���J4xʆ��/P�p�@�t퐄(��ī�o�D2BC��5��Yk"1/���%	v3�t�  ",�ri�y�!�3]o��in�m��+�q��.����:C�-�䉢��S����j�}�I�3A�)Oq�,�S����Z�>)�ϳpJ1���مn�����-��S�<Ԣ��a�\�����Ş4=�����\{F˯�+)��KI�J�ځ�{�OF8<z,Ҽ&EfVNN�0|]<w:�x�]�V��;���Ӧ���\|Z��0[����	��cݍ�u����S�|JY%T��BPe.��xu	���S8�/ #O�)R�^Ƒ����"X��[��Q[R�7�� ߌ���E����F7G#+�Ǘ0z�cULjaGkƊ~F˯�+)�"j���b7|#9���|�au�(Z��I�V�~��TD���rs�i���`�M�	=̞��>���ԜF����am�Za(􆿳�ټ*w2�56E[��\ �����^��]���>����C����N4������[�]�!����M[��Ǣk/�z�xEQv�ј�"��Z鎬�����X���*�Lt�2�t��|g�Y�'���Xw�E�i�m}6	��	Mk�rc��Et������2�~�7���e:[e��m=j��S
���t�  ",�������Ls�F�%ܪ���PL~΄gO�3f��*����"�Q:�{�1��9�����u�A��c�@�F�V�5����`K�aVD�C��l"�u<�rם4�S��ł�!r��Z����p��]|��L�o氶�#7�hY����r��4V�H�%ht[����}����g������(���B���ި���pj2�q�*t�ܶW�k (���B��ɓ�~Ҡ	u{ᵿ����0yI��j�Ib����rs�i�jf� l�Ǜ������CyW�f�tR�wX��}�
�?�k {P@2���4��)�ep�G;w�b!��uፍkv޶Gl7�|g�)���U,�(�)8���0y�	�C�u)�6�3A�)OqЈ�&��g3�g��U-�e,%�0g����ʐ��$���Z��o|VO�⅘�P"G�wk�١��	;q��^̽1��R��ӟ-�F`���G���`y����@����gG�C�cC݌1�"���y��Fp����f���,(���B���ި����x�3�Aga(􆿳���2����.���;��\u-/���yF��6�xZ��j�
�iB{�Z�_��㶢�&-���x�F`���G���`y���h}Nw��諚��y�[�!�TC��\[$Q��
�̞��>���ԜF��g.�~R���w�K�})9ͬ果�k�V\ިg��U-�e,%�0g����Ed��>�^u��v��=��b�Bϱ���w�K����+��dЧ^{�j�~m*�S%�,6KX�#���x.�Knq'��������d�a�4$�b!��u፸�Aݡ���Ƽ4g�'���Xw���,D���Uo�B��+ H�d�٣���N N�S��t��������ʓ���=�^�)�ό���.Ӈȓ�iӚ/`� �EJ�:��S*�IX0F�MV�ҁGG�.Mm-;�d�G}%����3f)-��^8 TŗF&�.S���"sS<�0�zG����ZAL�:!�`�(i3���y��lD�	Sz��
�GBQQY����#H�Yg�yi��v��BPlLO+�#}�{��7�i'�A
��ih�\�my$�N��o�/���;��(1l�jG���Z��o�̟�1dN�<@Iv��nt=:��:5A��p��;�/s�1��pn��>�my$�N��o�/���;���>]&���F�x��&����瑃�dN�<@Iv��nt=:��:5A��p�x���y!�`�(i3k������8���[{/;k+Q�h'�Ȝx�5W ��̫(�8�u?��I���?B��#Ɵe�*|�÷�Wе ;�jmT�#��"����G��Hb� h�ҩ�X19�-.|}�íN=]a��o���T/Pr
�ҙ�� л��Ԇo�	���q�ӘS��H����hzg���l�
@\ٍ�I�Ūe߰�	���1tSjv�!�`�(i3��;��̟�1����* 2|�:�c��	>�������Ra])n#���r����,\ͨ܉p�T�8����lr�{��|e��0�U+�qbp@�!�`�(i3��Ě���ž_�F��H����hzg�����U�._��I�Ūe߰�	���1tSjv�!�`�(i3졾�8 &����j�����3A�)OqO�5���1tSjv�!�`�(i3|�au�(Z��M�Γ�va�r\���
�oz˸ם:�c��	>������
�:qEp'{w#/ B!�`�(i3��=m緒�!v�/FY�a�E�Rq���my$�N��o�/���;!�`�(i3$f��_Ub�F�S�1 �fĉ>99��j���Gp!�`�(i3�2��Ȅ&N.Q�NJ�zQ!�`�(i3졾�8 &F;p�	l�
@\م�ԜF��}�����Hٚ�-����!�`�(i3��=m緒Sr��3�r\�����p��b���ez8�US�6 y2��R�՝� s�#���k$ �B�'��a���p��b���ez8�US�E�g�������(ӈ���m�r����
�:qEp:䩒=]'!�`�(i3��5��(���Z��o�XƤ5_���>�4No)�T*�c���-/a8!�`�(i3�3�7d`yu-/���y���!^��7���өzW�&��F�u��r��!�`�(i3rI�F����ez8�US��o�k��e�@�m�W#����#�=3!�`�(i3�����!�`�(i3���>]&���F�x��&�lr�{��|e��0�U+�qbp@�!�`�(i3HN��R��bP�63Z�t���%>�rG�@�	����!�`�(i31u_������]v_��,��q͛�����X�����a�ݚ�Н�|D
�W�ɪ
�oz˸�1�"���*8j��4	���_�239@��C2K���l��#��I�XƤ5_���Q����ݗAn�W��B� �b��!�`�(i3?�� Y��v�8�UG�����ݚ�Н�$f��_Ub����pT�HN��R��F F�E̠$f��_Ub����pT��5ߧE4��\E�W��4b��Q+��
�J�*���z臋�Ϝp��'\��i�x���y�p������!v�/FY�j]z�D;�*j2⎜@��'\��i�`8zo8�ǻOC�]@\��p��b���ez8�US�}o���,Ҫe���;�$븍���&|�2#<>�IX0F�MV-T������èV�5�5���/9�=eSe.��a��o���H�RtV�^L�J)���� \LÐI�q����`���*1?V��j�cI�ۯQ=�s?߫J��5���J>n���e�S�[�;.Z��ܽ��}Dq�f��\!�U��0�|�_�mS8<�n�ݚ�Н��tSk�N����C.�u`oPϞX�o|3��b�Bϱ�j�n�y�1�>`�nT:��g�XWfĉ>99��A0ok��$f��_Ub��7��G_���;�P�t�5�׹�8@CHU��!7D�I@O@ТKH�{?��j.;]'\gWg��	�Z�kfc�?)zni��`���φ��<�6��pɒu����Wa����'ž1�|�'����z.��W��!�`�(i3����j��3���B[=����e���A��s�R�b>3��g�d�tu��B<�D-���$�\%e��}Dq�f������AI��Uo��ƍ2���lī�=m緒X�X�pF�{_8�Y��=�}�Vݨ!��"� +}0�ʂ�j�Ï��	�l�lM�3 zM#��m����F�P�7��S��h��d\��H����o�γ�ha��o���H�RtV�^��=m緒X�X�pF�]�!��	Ǹ�y85������Sr��3E�¸>`!;�jmT�#�2��G��!v�/FY��Ei�g.գg��L�*���/r��X��|~����7�i'�f���Q5�Z���#�H�Ћ�r�H�RtV�^vx��c6���J����n��뾦�!�`�(i3�5ߧE4��!�`�(i3�v{A,�*��9_s�v�a��o���H�RtV�^>�Q�c6��xp�"�/ܲ�ۗ�DC�	��uc$f��_Ub�F�S�1 �t�td���5��Ě����E�i�m}6O�D mWN��ܐ�}ī��K��M����[*�q�K���g=-C ��U�