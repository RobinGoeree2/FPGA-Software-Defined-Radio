��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����⽸���D��6T�8�{N�/i�kf�!�6��̋"X��:�����\N(h�-����}!���1�����4�0���S��k��Xd�d���{�8�%���AHǚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
|)t�]з;�Y7�^(Q�`QԤq(�"1d��_��M�oЧu�Dt�2�3z����.�`�9��8I����w�义=� ��%��3�<w�ce'�j�A3N ��>Q_�1*�ǜ���*��'�G�BL^�#(��xw���ʉ�T sV_UC���9RC-^Rǽ��;�E>�h/3E7�p��K���F/m��:|�FK�l:p��ZvH�YC��c�a �~���E�O�5nʭWv�,�����?oB��h2�UЩ�*�yr��8\�`K��l��p?�WK�t`��bis�� ��9��O̢~�x�W�s;��4�l�Ȱ�g)�"�2�^���v-�YYB�Uӣ�Ԉ%H���f�P���n|��Ł��#���	d.������o	z���P�׻{��ӟ��48���-.��S��d���#�Vm�_F� �7`����SODt>)_�ZT�&�S�g�I:YS��s�] �ýW`G�I��Ow0z�B�w 4k��B�@7�|4��5.�(o�MT2	؟/�O�9�y��h�\���v�+]8b�u��n�����C����f�2�����V�KG��2�xc�i����n��WvK&�;���-.(��|A1�%�ی)�nu�
�3NN;C�,��(?yR�b��~�wP���'����������5h�^o�aS/��I^7]�~�p)@w�5hZ�'�{��6?�  '�f�U�7=��[���1�'Z�"��h�Ԓ��\��}U�2��d��0b�~��k�}�m��&�^���X���Z�A+�]`ۄBV�l,�+_?��Z�G��>}Ga�(�m�LD=}&�yc���	S�P�����OxZ�y��cD6��e���Y�?��g.�'�2�C>�@��j��>�dH�H�/�N�(e�5΅��8���	�?v2�+�{-]�>��м�oe����������vɌVJ�A�Ԫ��C�r�.�E���>$D͵y�:�VOf�ȋK��z(�3E�9�1��FS�����ث#YSs���'4Mϑnm�Yhஆaf$��D��H�" �����)`��D�Ѧ��AK�y��5�1�N"T S��%iK���|��W@_�E(�"���eq��L����1`��z�/��Xq�`n�����mp�9�`Jm� ��b��AKBV&P��">�gp�q���x�߮β��"�E��-�JC��0�x˫�Ka+�N��֣S]�4���%c��~}�5G����e�Mt����39���8�oY�����6,Cq''y�=Zi�0�{VX����y��ABߡ����K��4һV�!�G�J.���.�����v�g�D�gy��"�_�`.�"YvXM�ռbs������_��4�"œ`t諁nd�A2��j�5Zʐ�j�K=��I+�e�t��A��h�7jnD P��#��7�#s����d����<��;o@�-g~��E�f��q�2(��"%�R^8�J�:��T:��@F������k��2+%M;�`����U�t&�MnnrW>bU�{l#aY��J��&Gh�J`����^���ݲ���~y-��sj��Mz�s�W��^AD�?��sԯ��Ŝ�9����@��} 5y�7ZJg�n��j`�0�PKK�Y\�)��NX�*����D���F&��p
�v]s��
��N'��1�{�0�J!��dYU�wJ�Ze���7gh��;p~�� F����Z(K>|wy]�?�.&}�M����w�}c��R*Lq��%NP�:q�;��X[M���Gր (5Ez̀�^�6��ī�?{a7���֧,}���K�)�u�KW��&؏&�i�p9���$]�amu�AQ�\��83�ӡ��mEh��4a$�w��Is\�:��C�$��#�9�X�5+zy.�J��&
mt=�/���R��S?Y��{��0:^ �q�p������]u�P����ۡ�Jxm���XeY�C r,�m1�'�H�Z��Ld1�.�tp{�FKQ���������vYKb5ȩ`t��gAu����c)��s�c|���W�.��	����1�{���vr���ҍ����;;��ϱb^51R�k�!nU��,?������l�{k��_�
S]�:���Br_���Xg�?�a��!���*=KQM�����I�}�9Hj+x<�����;2�Pb���Tm�C+���./�ts��l��Bs�!�HOP[����QN�7h��+1Rƈ�c��a��/.5���9���ʇTW�-җ��u�7��{�ɍ=��J�^}^�5_Yʊ�b���	A҉������Pr6M^YEe9D�_��G7}�#�hT����^pv��ڶb�	�}1�ɘXe��[�%�eh��䃴�\�q��,3?Cג��t��0��\�tD�K��| f�9�H<(�0Ы`�|H�d��!�f��.܈��o	A]�qL`�/}��Ff�1�|���%�;�� ���-#��2��y~���kq��6FKl����`������E&}H��?��g�Ճ*@sq�K�����@��9D�i;����).7�iX���0���M�Wse���(��ݵl~wva���}�Rs�8/�7$O��gE�f3��$vC"����=���;��P2Յ\-"����QKM+� �ːs���s��6T��c5>�o��z����q@�,	���?c|\SܿǦ1]��LJ.�ܪ;�ך���^9����!� K3���i��g�-�wW�+�Q�u���=h{P�3�k8������iT��ٳ~=��Y��H�n/o>X��'`r���q��� �������n�Kՠ0��#�j����c&�����F�[`|G �����İ/�7����N�Q�N�΢Ĕ�&��TCC��.x���V�<�8t�t�����r�	;�|W�a�L��[G|+��z�?��Qp$��T&ihC�vx�CІ��H�����,���뫧]�k����Ϙ�{�F	
$�����j�Fy�dF_��b���T��8�: �|�v��TX�~����u@���=,C�셹q�tOHnT�=�J��Sq2n���U�������
"k~_w'�3�F��J�։�r��oύ�ǳo!�j)��Q^H���i	m��tU	᠀�BPz��l��s  c!�a.9��_�S�Y�=��N=?���2c�R�;�㯧�~@ې�$T���O΁jڸӣ����qy_J�V�\6C
�}�|�,����j�FJQ�Ӗ5�D�-�ң?�:W_7��I~).��q�Q����\L'?0����r~9�Cs�OG4!seӚ�����.�H�j7�^�p��4���	LV���38Zy�"��w$I��O���s�T�c������/��\�1�o6����4Dl@'P���z�Piհ�8=*� ���%N}�m�Um)Ǒ�pEߠ�	z���˯���aL~S�P�]��i�A��{#��f��<d�T�qlu0�˗�ʋ#���L;���RG�D%���_봺&�]�=
+�Ɨ��UϷ��d݀,���E��fK9�jaL߈-��;�x���!���'GhCg1DW4��a���,Kb��9%��4VQYS�����p
�E�@@�&+wbJ�sG����Y^%G ^�\���j�.ljUD�}�����52�k�t_$�$�6CmWi�Qa1�[}X�d�'+o-����k��� ��Kc��;*_����붉X�~��;g�)���CÚ_�{��ňw�m��;��+���j�v�?d;h��_�]��bMɕ�P�+}Kq�Ӗ�Q� ���}�Rd��<Ct�oZ�$ù��$2ܒ�0(�UE3JP�A�	Q8�����,����ȸ���Ґ��L�g����~�"H�tv#��ltB���qdMɪ	:`\� ��l�	�P��Զ��1"D�a�k�#��� (�Q�Y�,IH�o�'�P� AP��q�l���AHvľ�ќ/%��Q��A��V(!��9��f=�X_�%̛���`� ��1
G�Ai���9��(����<�0��f��� �����]�6��G��K;u����q��;(���͍�p��OlFo�q��V���m�I�IӓY��0\1?�{/Կ \YUms��7�$-Iq�A��x+x���[�7f5i*�����:ƭ@}���:Q���T{^	�ꦑ��x�����L!9���!��8����j(��0�~s�t�
��A⵨�Ȉ��9�|i'����F>�s�n��	#p��e ̀O[Sl�z��I6؜j���UUo ����Ш\E�����x�n��P��š����b�"�K"_ ߤ:�^�SS(��0���C�^�,\�_)S`���L�99J��A�F�d:�u��ТA�3c��G�������[�3��q��g�#߬Ŀ���|�7�J=4?Y@�zA&�p�h~ap�`\M�0�nҐ������I��|��L#gU�k�˄}�,L v.��.�Q�A��D�Y��rYp�P>������WA[m.n���z�p��>��EQ-�CM�	b��y��FZ4Ŀ}1k���©(��F�-��^,�>[���P�/�������^�����Ux�غw蹵u`_G0��dכ5��屙��l暠6��n�|\�[/ɨ
�fy�����*S ��~���Er~	
�9�#7`͔�-v;�p3�6l,&�u��1���_���i�)�~�:���j^.Ѻ�e�A�z0�����e��7.�l5��P�!ä�}0��x�Ȩ_s�m�5
gζ+jK���\�K~��C�(�Xϯ�O]�e��v�d����%� �������C��Ѡ^����&�WL��K92sOt8-)l���;_�ׁn�î��$��9�$� �?ewWܟ������u���7tVͶ��dfv�����t ���4���#[�q��7]Q��V`�*[�Сͤ���z�3�F�z���]�K %���ʲN����=hIqf�V7��,��`���mM2	$]�b�<�d���3�4���nJ���:��h�����y ����"2����L����.�?9{�*^T�Ôg���7Ղ[��g��5C�E2�[܋3���h��L���*aB<7h�\y:.�!� _�(�Q.��#߯��ϡA\ K�̒׎x�p� �G`������;\f7�s�b��$s�m20`p�#n����z��B$��Ěϓ,E��4A�c�W�O�n�}�jj������V��?�r�@�Ȩѹ-���,�K��U+���l�Y7
��A�B*��>���螥3�@�>V����,��8�hB}!�4���pD}�9�N����g*&���H���,F[�b�$ڣ+�@�k��|�*-ڐ� tڕ�e)Fۜʖ�߬��b�]9���'�␆�5�2~}j�� ^��+Nv�ܬ��OH�E��|�Eٯ�˖��C��k�ˣge�w�v
א���ϊ��qeb��L(�n����\�u��aU���.k����/I� m�t�2�9������	��4���qW�C!��I�[WT=�v������@�E..��ޜ6ɂq�I*��U�U��P��Vz�]�,�t�9&��]Dw��3����@��Tv1���d�� ���xԨ��pv��p֬S5:+yO��3ۇ����n=�-p��nϘ�1��A|�z��Mv�7�nᕺ��N*n�0F�ȊN T����|;%R�����D���8O���&�B�벁7FCHq]dH쁣��:ZGм���\��\�h��5���w��e�Hɔ�9}���Tk V�m����z��@`���E,�̞=!��;h�����y"�ёx� h$����2��Z.z��.J���Jk�-m����aHyg��sz���)���[�W�v~(����G''�8C�G>%�آ��rļg�ܭ�G���GS_����;|�Z���%��U�,�؉��Z��3�l7_�bA�j��y����Z����\������d|"w'��BfP�T�N_���oM�ӫ��q����v���sdf�s��p��S�H���	�m�?� �IF@�[�$��׼��T�}sz-_�4�E�0E�iq����G7��}��9��A����C5�Q����g9�n1=9g�,�a�WQ�j������(NEA�ޤ�Ed	�ȑ�b�#3���Z��6�d���e�k���=��~,˔�,T�/��$9����ב������×y�2�Ŵ�2�F��~p|k�Krw�������owb|g>ֲ��$�j��s��6�*�UO��PȍU�������i��ܿ<��7�u32��t�#!8M�i��f�t�AT�P���~
��� 2��3�k.��}��N�����f��4<�����w�u����T�U��z��E�ճ�:м�?h���p6ȅ�4*��Q�3dB���W��hͿ����	qw��W��9���:,[Ok?��3y�,�ᬺ���p�5�&n���K���������siCO��kk�(Q�3�[��*x��-[*Z�!�����Ĕ��o�m�Qe��2�o &>k�K�Ѯs��L�~��T����>�\����ɟ�jC�.	$����m��2[����fN�!�q�媕=��t΂�7%9�V��#�We��!���F鈀���A��܆ȧ�0PZ�ΤSc�"������~ щ�İ������*�/9y�2�Ř"�1���q����U�B����4�%�Y��>�)�&|y��<�J�C�։��,X~���	E���·ځ�}������)��O�;Z�47�W76�XW��P�U����\<�ycyȶ�P ׄ��/τ���������@e8�(҉c>h�Mg�)�+�6�l������d��f�J��x�[�9�Oo��ԡ���PoP��gf���E��Z	"*��כ�E_ee�������¡��u�p,P�i���_'���I�l�j��	���`6&W&���J�uş����5�z�t�|I�;��aTm+��j�~�ی��z�g�<P�h��5���Z.��*�΀�I*��m���}#����l-Lu��X`q��L�*�$���������P����c��i���^���4a�PF��;H{,P�0^�礦J�A&��Ʉ�Հt��y�v�i������OP�D�����be���%O�Y��qf} ��O���Ж�CG������P�9D��t���1��y~)�<�nfذU�= ӳ��\�Hh��
���m^���A��:r���:n{J�eZ��t�nasA��zm��!G�A8�~�`59��f�B{���G6��Tvglh��6#*�.٢(�)Z$�&'az%�O�(f~5���pL
˗rn7�M+q��d4�� �$�g���8�{DQ�hS�+@�3��Ф+k|LZT�B�Q��T�!��Vi��#S"<1f�~��s�?s>���T��F�a�
/>��5>)-�;�:��u.·�tӦ�.���/T���3��J-d|'~O�����n��ݣ�V�F�k����W �C@�
�2x�C%�����;j�@���/6gx��<����Oĩ������p�T&�1���������ېER��^�`��^�W���L�PNB� ���fˣ��'�.�@�j\�i>'h��+�<,���B��� HqM�M�(MU�f���9��p�+���~B<L��Ů�y��ժ���"س��RT~��^l���C����3[�lKPM�Âb�i�l���i�H���I�IЊzf����->$X��BE$�ƙ�U�P�e��z�����0M(�JAK�qx���'J�QU�ҽ�%��ۓ�ܧ
>�3�0�O��	
��{�ЈW��p�:���Z7��OHZ��/nv�2�]'��I}�1�!�.Э����|���|$(������HE����;�s�]���H�ߠm�>w����B ��Cl�_�������ঀBڂ,'G��n����C��aC���AJ3�B�g3�[-/��=� �o0��n�d�sh�U�F��C�M�NSN�H�~������2S
���/�̫�l����E�8�Ӿ��j���E��d�;�����+6e�KH	X�7p�q�?�W$V{dl�(��y�[Αg9����@3QE�ae/�
r6����G�gw���ݰ`*��ɒC�Ȗ�	�m!.t�x��vn��b2�o�[�|��t|����8�Y��G2t�q��a��0�&*[�`O)�ȯ�O��֊����%[�4��)Ηji4"�-rr�ڕd�&��MS(��WӁ<����n���- '����H�1bχ���q#!8�'�`p%��
�Wv���%�Cs����=Q��M��}�\`O|󔂮��*���/�ڹZ�n�����!��o˱��5I�Y��������_n �"�|lu��Дa	�;��z��Ɂ��"�`���Z�su~� o����$�*P���{s�.�w���`"k��>�͚�l�	�-k�`2Ų_9ޛ�\י��.�'�ǁ�"s�/����Ȉ����pqG3��	�5��r�(��	�����A�f������I�c:�3ȟ�k��0�\��]��"{hP�2J�w�G��/)�D�`ƫ��܎蘆4z���� 3ZI�&(�4�-m��C���=_���<'�����{��'W��lk-�P����(�҇?�mmR3I��M������9��Ќ�t�=���B$xf7�3���&&�S}"�B����_q�j �ߖ�xozc�n�+{�&%�!ʇ�yD�#��#�����u����o�d��zy-K�WԖ�%�"I��K!ڣ���Rt�JkutV�	�?q�Yw���/Y��"R�!L����?K��ˍ��k�]�i� �K,\цl�-�l�@_$B���OK蕓��S
y��>�Rӄ�B���>�Q�n���#R�gFb����G\�hyn�}�;��f�A�n��pC���8�d*S��-�=>m�kp����H2��IZ)I�<-�ҥ�VJ�����p�^g�<�G9�y�4<�fz�yb�;�jl�r�,�s�#��1k�����GM8�F1{����M��<�SE��W��F�[�QL�L1BVߤ
��N������<z�9hW`3��B��\לM�W�L�wdDE�F�]���»8��&�y-��]��~������2ߨ�s5����	�S�Td��1�E�1�.�E&���5�
�5w�[�tO.A��⽤Ӽ������h6Bp_�>a�g8qd��z��oa�.���l�����y��y�q��\lP�_r�D��Y�����y��x,OC��M���u���+d��y.q��ρ4� ��������#V�ʕ�9I4�>����T��d]������o���<���]c-K5Qy�Ĥ�#ʶ] �C��T�2�K?<�a�+��'�WE�~ٹex��od6MO����W�����j�����97������b�e�	�e�82
>D� $��={�z�Sd>-/#�Y�Ʀ�lM[�!�5"6ِ�n�� ���0�Dju�䘕O�G)h�Ƌ0c4�΍nyX��dКt���$ND�j��N��2*J�<��X$Vu���7��pdl$=ylI
���F}�S7{���︪O̏�_.>�y�R
�.Z}�N��
A����O�T���H�%�e%�����`�n:%�h�)��g8kn؝���/m��X�%�_���A�2˰�����7�q_H����'�#K�G��Ł��}-�r�[4����~�4�K�'3��,�Җ�FK˚�\򖝕d2J�E�u�������c���i��Ї-���Va�W	��i�a�T"�6T�v��5��3:��pYX�VxK �
�i�Qc}��_��5�V�X�f�Zu1rW�>�{�|t�D}�_��^dhfp`{'�����m���cq�<���K��q�$��(��X�����p�oe�e5��vP�TQ1�Q2�pq��v�d�B��}�r����������'p<�_����=Rj9.��1r[��ܜ=-5��y��':�x"�����Ӷ[���fz��mY���2b0�ùc�ThRf�"�3E6���*O�-�
^����ʛ?"/��	H�t5�(d'u4OJ�+]�e�����r⍄���zu1R��A�zc� �L�2{V���r���O�B��|ftZ�̡�LmJ�ԡ�."矀�M/�$ �7O�@�C�D�9i�/L d[␆��.�\J-�W!��i�&g��u��&a�}��ʼ�o���1�wK��B�E��j�Ż$�ߋ�`�@$�3KR@r�܏���2�∴ 1="lA$����:�p���<�gK���Hr�,�3^J�v�~4��Y��bT+��|���a|?�U�c��ϯ@T�3Gf]B�6��=���D��x�Y��^|�E�A��W���fv�����c���@�6�m@AN-�KEU�Tv?��D�xswRPƽ�"�~�(v��o�Oh^ }����� :B\ا�p���m6�U`��P��R��b�����K�?u����h���z��i�)�;٠�LDJ���ș�	�	�Aa9[�?��
��ȕ��2N_�hh��L�ʪi��p,0��k�"ە0ʋ��r������	o-Fp���uC&K��~Y��|mRg��~�����{�*7��:{4�&���І���;����#����VE�B�[����t���U�|�Ҏ��ClUOt�_4�^���+�T%��(#~/������IJ}q�ht8/�!�]�{h:��+���=M��OV�M��,������J����F4�w��Et�� YLG��oyN�G3�Cö�d6.���� �O�ڋwG��?�4fP��$v�H<�OD2�����9F,w
\�BAsl�h��bjcKƈ_Dm���)���7镱�<�v�3��0><߮M�>x5r(4�+b&�f�1�2H�9�+X�\���h#�M_w@9;�_2� �u|��.�3�8����5�a������.���)f�lm�0^\n\e���)	x��@h�U����Uo��G/4��!�{TH}k+�=��)�z/ 7���B�}���l�7�v�@HG���\s+�Q+^�������M������������j�k��C�X��X-�ǭ����J�2�T��U��J-����� \դ�V�����%���ce��*�s����7�p��zl^ra�a܇y�!?E+%�//������ߙ|0�����7SX,%��^���\f�E���rǡ{ρ�5������i��,���Kge���pȚ�֩�5��-�x��'��eZ��n�Qa:U>^jпǱĽL�1
_��ɏ{�g�
+�-�'�D����ͺ�%h�Y�2�a��'�>�*���\^y����lC5]L�l��+Y
/�[E$��eYu��fx��ڸP�����_6'a�1\t�&|��7j�h���ҦiT�]|,T|2kQ?�a�W�UF܋�q�q��\`�Q$.���r�ʓ�*2�|Ûyi�݀��#�ǹ?ba���vHg��D{�6�J���]f��Z{`����$�8�����B�������z�\����K(sS$���4&,7���������+�H����A(�r��q/HN��}��x&t�T��C��q�^�sM��֊ǫ+Ǿ�^��4�Є/��^b�K]fa��vډ:,RZ%_L�"WgE���^����;-۝��J�)H�v���`�!c�pl^�Da3�Vԩ�����8�(����{!4���s�<+A��4�8?􋅽JO�tL�Z���Q�S`k[���}���	i��;�.��?e9��x����vv��g��n: z�˹���p�5֛��N�^f!��X�kR�@U�'�`#!@!�vg:��s�R�lꭕ�;Đ���A��G�4��X����3���r�r���k��|e*������؞���4A{H���<�-�L�Oԗ�3�ל�4[���Jُ/b���!8��^���
�6���T)�;¨��+�R$�Z�t�RrR�s�?g��H[ݸM,F�:���V%��hW����&l�_�c-�J%X�|��|�hja��E�{����9���/�4�B"�$7���x�"�R�@䂎`��gS3�[�����ͱk��$İV�Y��;kt��\VCs�NQ����C��W�� ��gM�}����A%�f���rO2�h+�֝�W�����L���ш����R��6J���@ʟoV�M��YQikK+����_�j���3l��=>�s�t��Y��0�� V�cf��A4%�eF)����o��ى����zeC�5��`mk:82Rg�_8�Q��Rb6�b�q(w�F����Xed�dS@(�u�P���Նq��G��׽�u�)*N����dqxb��z�$SfÜEҺ@{�M��G����`)+ЏOv&pd�lO�8{��/�Qj]��\HJ�=n��,`Q���g������i����P�ؕ�NT�D w8�`�uz���Z����f����ݑ�����QV�,��;��6�	E&���k0��Rd�%��>�%�#.��C���娧�5�(=�3�.���>�:Hb�@��ւt�����=�!+�x�h�^��V�[�3��
�1��:A9���������{~Y-�za����C�!~����)�TT��ʄ�li�ٔ�	�Fxp�:�ҋ�p큠�b01�g��ز�� �Z�e_��*�@#W)Uw��@!�q�G�;�-�#����*�RQ�VF������������Ѐ�:3�d�SECQ��&�\��*\�~����� zw���U�M%��W���:
Kj���e���Y�"x��dW�ǻ���6m��� w��>����FykV�o�u<vL��S ��W�#	��n��> V�����ǯQ��O���zp	�i�3�r�~�Ъ�׷�jXi�**@�H��Q�z ���&!,L�nWƝ@V�bK�#t��(���2S�˅���uJ�����c�5�={Y����L�^�7?���(������V�D���{p���A]� GKTI�����o/���&_��Ge�i�`Vc�ST��u�굯��v�m�_-��e�)�H�Oh5cw��lE:�,c� 2$��6�W{x�/�����X��.�19��(Mۄt��V�~b�B�l�sև�i\!��OF@+����lI2�	S���������9������z{]�҆���`�� Yf�3{]�EՔWȩ���}�@}��i7��̧7lH,E�N��Ѕ2�G��-g�˙����ܼŏۧ�ś��I��t�^Ϩ%R�.dĮ���h��I�
+��fr�#2u���nV�)91��w��Q@;&�/~{O��"Z5Dv@$�ds-��6�[FL���������O�~~J����=�H���촉ˈ#D�vb#O�xk��L"����1�!�IΦ�:��w+`�����;M|�ࡏvFg�}�ku�E��CH��g�?�s8b;Pz���������C跢����\��N2]�on���e���,SwS�#J�6I��p$PA.���7ۚ&N�r������Q�� �X�5��K�`��x��bOc�o_�SvWa�*���튈 #�]���7���ͩM:��ˇ�ıw?H���:��U,3���{�;Z� -�0[Xw�Ay?A����N�&X����~^m�w������xѵ�J��M��R�&an�y��r��7S,�ٝZ{������hԋ��񴎁3�.Nj_���q�������Ja����tQ����Ǿ�a�� I�ʍ�Nd���j/!OK�����G*(ω�g"ws��ڟ��;�;dg98�(R�3I�e��z$�^�Ra�kd�U�]g`	��gZ��-T|'���(�*<��8�s�͆�{pR��f��Be�n3���sO����%�������I+����[��17��9zV���V&��*��f .�G�x��O~�"�сaq��[t����Y>����OEQ%AIe�ݕy��HR�x��~Fʕ��w&z�ҵ��m_\�!v����vFue���s�:��$�fp�U�ϐ�����5�h�ڑ���B�{"���$���US_qt���a'��6a�r���`���k�A�O�P���P�w&t����!��.]d�j�i�Ll^XY7��)���p��f�<)9�����nW~Hk�O�����+��V���O����y���xms�ʶ�>��e�wl葪,���Z&�0wQF�&��oQ�=x�!���6`
��e{l�ȨX�Ǖϴ���`^�^;`Er�~��9�=�OV�5g9 b5u���F��ȹ���$�(*~��� a3��X��^��!�,V�b�1�iՎ�����T��$
9ED-��oJf_X�|p����Y��7*�<�w���).�4u�9a��Z��`�b��/��J[��Ob�9-%G���őb�^����1d�瀪�q\Fp��7V��Y��������+I�/�ν�_�I���N�ڛu�wpdx	N���-����S��b��f���,�,Y��Z@�g�C��������Dw�V��x�o503�S��zͶ���v]#{M��LS�����O�����F��1�6��)�T��G
�+3f�J�����p��;���*�yZ0�E���/�9"2��UFp��u6���`��Pn�mP�����݉��HVV��m;��*��9�A�n�Ɩ�9�� ��n��Æ$�=Ev�ۼfn��%Y-c��a��JY,w�`3�8�m�ƒ�r���C;Ek7K���$�]�g��k%"��Q�1���ȭ�> �v�����.�̜�`��Ar������&��sJ�����B�(N�������Zٕ�S�ّ@�DT��s�t���1��[��܋ �k��yȶ��%�a%���xi�|]����G���$���C:��� �Y~UG���5�|V�V��F1�l��6>���r
Խ�N��hp��ia�zk�da��s;�-*����t$�.���E�̓��pN5��W�*_""u��,�8�$�^$����'�u�>�t�}��.�B���Xa�O�b��7KOvm*kr�l�����a�Ndw�OvsB����؏;H����KC�5�4.\�h�`��I���+��aoa�:�J7�Y삢w��QߍԂ��af��%i�2FYnMO�^{s`)9��HS�F�����n�x�Z��d��wP�:�*ԯ���껥�C�p'q��%��?T�N lQSn�S�� ��=D�;�2���JLݫ��?"�$���E��No .�)�&�A�4�\V0�髉k��gKPl[�9�`;a���?&'�1EZ�#��]���c7q��>=Kr�ʈpD������0en��)(����V�ڬ`�mϲ��ii�iv��G�	�!�d�G]��� ,��+8�3����3i⼒<�Ğ��0�����Y�H��&z)��kPAǃ������_�I`Jpt'��dm�l����2�j��=:y)��3s<:�F���v�l��Ӫ-1���Hk���kg�ا�)���~a�e ]�?d"����<�+^VGL���4s��x��^:�c'��Ղ��2��$W�YL���L_6v�G���x+;��	��K>d�ml1e�,��m릭����(��u|oL��U��o�w���7��Q�</�eZ��ݨ �)�}F�
����/��Lg6v*�bM3D��~��Ow�S��,�N�G�X��w{��2� iwz�­����g=��r�ۨP��!�Wt:�I1!O�0�b�ޔ����J����	�C����E߉- {(3�x�������ǩ�9󥾛	�5�̡q�\O���6c��S������騸�q���ń�<�@-�0n��v�Y*��3~�p�s��L��R�L�W�����w
�Z�_ǲ�J��BNx��J��!`��Ɋފ݄��.�&U��R1}c�6]1��y/$H��hWN�բ�o��f�U<s���6��[$E����,֝-+�E��q������p5>���jQn91�����v.�d��X��8��;��>�}�v��#F�X���aݹl��V��ډ^Fʈ��Z=�����7�T;��L���s3�EE,��t���ȡE�F��%�Ǝ�!N����	R�JVg����}T���2+��
�ƽߡY򣭦+��R/�q�)Z�k�Au��Y�x���uS���sÝ�%2L�^Y�������I7�_-�@ң(�s�/� 1���#݂	Ls�2{��Ќbs��l4*8K�K���3��#���U��ک�[}�?)[(��d��6�.e���Wj��d4�+���r��J}��#�d�>�.t1H<�g���3,����4�=�e�����X��]�[�T;C���h���*�{`��uw�ݓ#�'R�H��{�xP�:$����w[��X�E�Pƴ>TLΑ����W��C��j�q�5�MU&���)[IV�%�� }�����6cˊ05�i�����J�m��+����Oyo�63>7��~���8 �5$^��$&�_�(�C���|�l���]T��/�K�	�g�T�h��I�Q�L��?n�����X_�%,�>���d�O�E����!f��
�oVH�O�v��a�"Dx�KGM'�Pq���!��_��3��ݵ+z#$į?r|��8�Y̹�H�Y;N�K�A��M�+��M�.M*�B�M��ߵ�c�->c#�b��A����y�9���3�Z���� M��#~y�m���t(����n�a�<ȳjo�Hx���u�$-�̩k�.����3��'��<���g��L���T�Ue�_�42.���D��>�&���M�r��"�8��2� ���f&�V��	˓RK�mQ�v���?���N�����a�G�]���n]��!=�ֶd苰1�Vf3���;��4Mm!$����ݿf��z�n�K:�Gc3۳f����7M'Xeʔ5�E�N���<�.w�Q�]�6�!���m���ˀ�E*x�O�g�[q����-W�Ocϩ	�_][��sY�Y����qJ��F��V�<{�i"/�j?��C������J�^�n���jT��C[`�!�qq�үj����/����/ �bNR�L���o�ό_eu��^Fn���*x�V��#pXHHL��	x�ll9�i����� ��h�h��@@��ʤxI*{{�G��י=�'��g�1�^(�O����SIꡃ�����7q�=ka���d���7L���zb�:��_���`0T���6�==���֗����_�`4��O�)j%l�̉Y���Π�Á0K(QzA
��|����UH4y�w�,�� �V=+U��>OC�vc��/&*Ѧ�Z<8Z�Oo�_V�Zz�U�_-|�8��@�����; ���t]��]uYz\*ޮL�E�H3>"��og��0����K�cX�O��x�7�&H��:�X�o +>	�m|�]�vF�=y8I�y�������U%P��2kVtu���50�T#�^��#��g�E����)�f�W-�O���"�0>���
(|WԂ��Vv����QPjp9��%/4��,�y��1y��M��sh3A��ܾ �vSTr�ln��6;P�<��%�/��U�ۙo(p����b�O�1 >c.yN+�3��3��ݗ�a��#����G�p�,G<h?�"qf�=��D��Hx������py�H94��uPl_02���>ۅn��<H�S�!n�4��<�*׋���b��s�eW���tO_i�~vifaJ���h琂L�j�ľx�/F�k�#� ��1�W�y���W��1�:@�z�Щ'�	2E�����>�%Vj�d�ׯ�[)ݝ�u�W5[�+��b�r��3����*|�'��Fָ���X�4�X���v���뤫1rSIv�r}��(�veċ��6�M�=���Th���!�e�����_,b���]�K�3ue�G��L�:���� ���#�N�����͘Png�ݿ˥OB|tf�\-J(X�mg$����t�.�y����[�¤,��ͣ��,�=��ƣ�`�غ�b
ﾹ �=\��@i	����Y�8��S�d���3!��
o��(�nԋ��W�v"Vc]4sRU/�1}��?����O6���~��/r#����4��8�Z�Z�X]��U��a%x"�PD�N�9�2G�H���,���b�����l��9�����dҺ`9�����'�>S�Ӌ�	���s<�2PQ��BE�E��l�s�K&��U�p�>P�
�km�l�O����k֮��%��e�/l�f�K�/#P�����f�u}"_�w�dY�����f(��ȹ��y+���n����5
�˧ϱ��IY�����޳���	S{]��c�Q��@�K@�>,�\�w�!�E�3q�Rj�����ޞ����m,�F ��Q�?X
�$��[f��3�Q�^��!�n���p���� Գi������p���*����vk�}�{�W�*�T�&V	`��p8��%��Anc/w�6�/AdңZ$��R�iD���DQy��� �?f_�D���,�Ba�߬F.T!��헪���$K���Ŝ{��A��[k�_���Dͦۗ,nko~XL0K`	��K�I�L����%���Z��2��-�"@tr�	��`Q�
$�)�����J���cy��	F.�����@���1�2�4�~�"����4 �bx�;T4�z/s;����r�~
^ힸ�~�ܗ����/�!�`W�\��8�|��U����C!bk$j�8�����%�Y��Q�Ŭ?��X�T��1--zIK�	����R<Nh��f�����������#z}�b}���rT���8������[�	b(�)�ތV=��a�f�"�f��/��E�e�?ӓ��9E�Om���
Ѭ�d�^4��X�ʊ�;R���UŐ�G�t��a�d ���
�\���5�b��G�oU菑v��D<myX�w�Z�\ �$LK#v���,څjn6��j|*g(��%���[��4��P�����V�:���1���99F��?x��$4޿JFEp��\���ؠPs�}3fυzr2�ɾ�Y&�&����`���NJYȚJ��K���\�P��D'<�(K���hi�*`�HV�Sr#�ʰ��+��3h<�!�hmb�QH3���#��i��̭fߛ�L���[��p�۬{z��@�|����Pg�G�F��ihm�b�/TH�{%�[O��N0��t6ʫ7<8��?�0f���Z��%�N�y[�V�͞ q�c7��	��4�)W�І�إ)?��e�΍V��2�,щ�MUKy��
�L�JLY�P���k	rBA����v`e뺺?b%��̟H����Q��ɉ�ƞ�)���yʝ� �ɋ���P#�!0�gf����q���W�7IY��+\��D-�Ș��¢���>�~o��60�쩲F�UP��:�	���q�ۺ�������y,4�u]X�W��cU�U�h��}�����wu}m����X/��ܩ)��EZb���{��`ˁ��d��x���"�D����j���Ɇ�Y>����ag���,��"%A��h�h�J��1F��"���l�G��l�a�0�b<.���qqC�)�YR ��>�6�Y�0�?�b��:������ȃ�Sڬ��tk�a��ǂ��]�'���LC��:m�R����~���c?��@澣�L,����y��$���"L#[�ֽĺq+�+�ϼ�Y�F��	qh����~Η��:'��]SP��ە���w�-[r�Ba��h�W˨W�E�*W���*�ow��2K�-Rb�c/Y?������+�v�/�DX��ꖞ��uh���h���ʥ��aKb��	j ��\�P��������2�D=쒦��r��\�?t ~a�
��7���9�'����>�W��������.J���썜�9,[@ؙ�Y�WZL�,s��j;Js�+����'}�51G��a�:���b�U0?������h��| �����p׈ţJ���u���$�w2n/AJ���gz�c�)`�� ��r_�L�,W����،*Z"!~��f8-�����Xƫ��]��_�LX,�3�Ѯ�m�m�=��+7��3x�jkS�#�p�AZaQ0�_��"YF�G+p����<�Kǘ��'�SlƇm�L7"("tۉ�.���KW++�
�;�QKތ�-�c�/�V[�m	+�W�k������C�b��?��UVn�ͧ>E�+f.7�( �˂��� x<�������BsnH�aI=cz�J�˃@2/����8�����{�L�5��z�&��KH��mH����J��G\�?��N��6j���Ҷ��i���3:ܲ�xX�/��ZzB,dG�m��n0�������K94o�� ����*%�FY�Q�µq�C#ly�ͅ�7�|���)��������qk���R��%��3���?d����D}�B8) /��Y����=�q��򬡼�"��_��?�s�M&of.�-R ��{���YRa�֠$��>,Q���y8n�̤��˪���8Tz�T�$�P�>��O�p�uW