��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���G�H�ƻ	�"�iQ�����3�7Q��㼫F|�ݽ0��@h ���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω����	8���/P�p��]��;�Iώx�t���E�L#uc��WŬ�+�-ޗ(huUPy�����h���!�}�1�:�Ω����	8���/P�p��]��;�I�����)O��Ξ4�"�\�� ���K�O�{��
2�D�� ���Jc\֣�I��B���t��|U|�/֚m� �+d��.8%D.��n�P��<�!Q������Ś��
��H,7���ZXWL�sZ�	!w���� �bRw�����IL�+�{Dr[��:�\��~���"��y0��9�QH��������\҂�% B]�pE(���B��|����<*�(�)TQ$|e�Ny5�7\F���r��RL�a)3���ʉ���Vu�?*tb_Rƚ4�%W��=n�nI�7C��H�pc;}
>2�%1[br�O��C��0��$�>��w�|(G֓�*d;��w�>��S������kk����a<ʍ���n �P
� �AH�W���,� �b5z�箲����Q���Ŕ�ԝF@�4%���w�K�@p��:p�3�����v�/�ҥ{E�?��RL�a)ѻtUWR��]��5t��^���Y���t�&�7C��Hl�>7��yx_/�Z�s�	�=5�NUD60L�U<���;�e��e����[�/��2r�O��C��0���df���z�!%���`�򾄖�u���;�����6�b'1�}��)��gi�HF��eUٻo���mi��*	�ť�.^�i��' 1wH�x�xs��3�<A��z����
a�������~�+��,/,����W >g1�]l�&Y��F}갨y�����# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��`y��f2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�����g��~�X�x��S|�m����Y�{'%s#K�v]|nf<�,=K�F��N��j��D���s�촜g1��rN�.[4<�6��Mz�8A�P�](���࢜p���p��^2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>�ϜT��:�E�>�5�4W�g`%J��N�9��N�^#?���E:�J�k �?!R��	k�9ːh���%��A�뱛+ƯE1j$,�����������ӯ������@	�J��l-[�v:v��M�H
�}ʊI�٦�D�`F��al����Fv��ߑ9��E|+�5�(�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���i��'��'[J�pO����1V�[���BV�GI$��ǂcY�~�ː<��2OYTT \��{9�k*���開<u��R��0�z}�J�f4f*��x�]�V����<+���U��\�v�w�?�b�>��}�+�r1D��y���T�Ŭ��ؿ2�%��ĕT�u |�&��R�{tks蠗�ةO�ݏ��9)�PP5�q�*�҆%�t�1���Hػo�V��+~N�.[4<�6��Mz�8A�P�](��h &�=p
����L�]�b�֘m��+?��bV��ݚt�  ",��`&�`�y-2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���\��tT��kU�!�J��E	�]��c ����ǆ	p���Op�ե[��S`�^yLٌKp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ����"��yݞƼ�Fm��.v��x�]�V���G�a��-W`������a�"�Z�>)��hC$?���;���EWrg��w�-�W	�I]����2N��n�lN�Eï.O��EB��5F:	����n4s1�ЂDa��(�_�R�G޼QE1���E�x�u5�����}Y�8?�pu��<���Ŝ�����Uh1�[��(����#�a�Ą���ee��U`:,��H�RtV�^$ Hl�]��rE�W�xWQL&�v��H{�T�T��)Q��QL&�v��Hce'a� /k�V�O��|"�_`�CÕM�yx�,�Gz�7Jg��q{�).+�Ȝ"Cߚ9$f��_Ub��7��G_��Ct�w#��@������37y�����:��5f/��|��I�.�����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h��9��ӼN���,��o���&W,�mI�p�\q��+��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hN>�4�
��l��d��|)?����t}9"hǸC�Q�5}�m&��߁�1�b9���M��A���"�g��bc��[�Bf�^:/��T�n*�N}�m��{���-����c�8(;��P/;D����i����R��$�Qu��((w��|I�*S ��1Y�ΊS&!�`�(i3�R�Q���=�>0n����|0��.���Q�q �԰DH� ��b�FP&[J@&�4�b9���l�{:�1���$�Qu�&�<��G��d�ů��z��_#Ԡ�O5�E�i��K�� d=��¾ȼ��S�ș�֩Y�3-K7͍����	&��N�S,I0��ݨ_F���m¡�R'cf��_n�����a6#nk�u�+�v��Q?M8�f2`Y)hZe���i�z5��>��(��Z!�`�(i3K ���x�?�@E�w:Ԇ���� ���y2v�W�+3_�?���cn�:�U�z����ݨ_F���m¡�����z���:,c����vH�42��F���m¡��S�ș�֩Y�3-K7͍����	&��;b�-�2�'{w#/ B��S�ș&>K}8��.KH\���k�A�]�����}Dq�f��#^���,�Z��xu�T�?� ��}Dq�f��5ߧE4��HN��R���מu��� �H�0��
��X��rJ���M X>ݞƼ�Fm�[�?}õ=o E��h��^�R�@�6�֐����o���uRTV�ݵ��y�4r7�,Bp��S�\E�W��4b��S�����H�
B#��Mz�8A�P�](��h &�=p-�b�+�