��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���G�H�ƻ	�"�iQ�����3�7Q��㼫F|�ݽ0��@h ���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω� C�`N��D���ÿ0�^��p���Q� ���6��H4ي��2_)��:B!�b�ؐ:�{T�{df�r�<�XD�* O�:��9M��K�:R��,1E�I�?g�f��r�F�5��I^ξ��ݴg��S�ZC3�����U���T���딣0&_���X0���2|	p��rw@	@us���
���m�jm\J�ԭyq�`݊�|���"rG�
���}�\�.�DV	��dU�;�\��^�� ���K�}M^UQ�S��)�e
�9��Ax!P����,��*�b؏�@�~�S�`\��Yi?��n;�|-���g]����g�����fP����IL�+��ץ9�^kh�u��<��T��� �}+~�8Ó B]�pE(���B��|�(����5�?�J�Ń��ɖ�2i�螘c&��(�R4�K��9�ĒTC��0��$�>��w�����N%x�g�u���;�Թ!o�o,%H�%��1z�:맷3%�!Bd�&Z��K�s'Mm��+|sL'���oֲ󄰊f�'2,�
�Ɍb�a���q�©������5X�/x��-w}�~�����(�1�e+Q��k�8���҆�|n�����|Hj`�~^T�ɴ�5���g��J�Й�m�z\H�� 0��~����p�:�C��JS�Ȕ*Ĥf���J�D{g�P�r�|Aښt�  ",��9���1� c��(�U����	x]�<���e�P����>�]!�ՄN�Ӿ��)�$�����PГ��0�w&��EO�{�������E��sޜ��*�c�N!ͬ鏈wƠ��ѹ?�����qU�%��Sr�'hJ�.;��L�OT�+?3�l� c��(�U����	x]�����O���8�t	;N���=��B�3ʦU�:�%�+M��m}on���b='��\�4�sW c`k��TT	q��$f��Z��FUR�.�;�~�MUs �ˠ{�t!�.�r�c^�e���zǒBs�&���b�!���<< �sN۪�c�	u�~Rp�,k���%k�&ָ��sE��D�őⴔIꈸV�MT7xB2I�d�HnULkIh��:h
�[ϸ��W�A��S;CM���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�
+&�s�A�F�7���3�GXS����E@��~���($�J.���
�=W�֯��i@F�5�=h�GD�#�̔"v�lf)@̲#;���(�s�-���f�i\􁗊�n��\v;V[���b�/r���q P�^�&d�A|�1�:�Ω��]��
��rE���ƪ�(����D�I�?g�f{ì(Q[nS5H�j.F�6�Z��'i�tw:g+��T��٤�2[51g��f�PH2E���ƪϤ�Yk"1/��L�lW��+�va��2鍔�	g\A�Ny5��	g�y�+��T��٤�2[51g���i��T!ea�8���*���g S��/P�pݒW*g;X����ˉ�1�:�Ω� C�`N��D���ÿ0�^��p�����rYd�ea�;y� ����t����M��҇+:|8X����\�vňu�,�s�h�' L� U��֜��3�a�\����Ŵ�(??a,8֩]=$����N�a�A ��E+���XP���4֔ʽ�I7��-5eE(��o���&��J��Vǃ���^�F��M֋)�[���6JHn��z�ji�gw�<�6�Q=\K��OL��4��D@��Z�y�#^�h�S{�5��lW0�>���'hZ���溂�U~܎VV��EfVNN��F��F\4];ˍH�7��_��T*�7⌹I�;���[���wK35������8�TP:(�������aB7!0[����	��N�Ae�#��5?�&P-�^��Hm��e.��xu	�n�-�6��
�jW��D���M��ҹf�f3'���F���;�¬pX��g��U-�e�,���6+�+�uB;y��Yܘ@��@IE�U��n�-�6��
�jW��D���M��ҹf�f3'��$Ι��o;�¬pX��g��U-�eן�-�Q�Z�ǩGY<��z��}�\w��0]��0�&�ͭ�o��C!T*�q���U�&��GE<�N�By3��<Z鎬����y��|�!�ptӱ1R�m��+++�i'��Cx�"T4�^�o�M�<�/��욷NË�����8��z{��E�EYZ/�矘��-n��I�?g�f��r�F�5��I^ξ��ݴg��S�ZCR;�{m�B��Ҝ��a�N�}��t_���Յ;��n�a�x�a(􆿳��Ak�y�y/��=��K���c|�7����+��_�F�����CY���<�;�L���9��Xv7�j�i���TR�^Ƒ�ӽ�}^v��Z鎬�������(���`$�P.eE���lC��U�T�\ ��y�.�`L⯣�v[����_��ƕW��V�6IWJE�$��dg0J/��=��K�E��{#6�ae�ˑ���CY���<�I����"�ή.mH^�+��@}�M�U/��Dk�9�{u�݁.�qO�.= ���V�6IWJE�r���秹�3I^�v�%j���_E��V�F�r�f�t��6��	���`y�����g�,P�n�Ͱ��Le�2l��4�y��ɦ�@^7&ģM�'n�^0o�<:�W�_ĵn(���˧�0z�cULjaGkƊ~F˯�+)�"j���b7|#9���b!��u�^�9.�JQ�"�y���[�ͧ�?Y�f�kN�ı&l����[}�@��L}�
�?�$���]׽���'�e��`�)�	�%{�;����f�kN�ı&l����[}�@��L�@����gG��l��`�����C�#�,Z鎬�������(���P����ˮ��lC��U�T�\ ��i3�|)sՀ�T:���V�L-]�#Ka�	r�&B"K�͢'����&���Z02��`�z��GZ>.�02�0]�J�$��Xo��I;��?�;���[���Ki0j@$��U� ���_;���[���(��$������l��p8�Kj��#�M��	GT)y�h��=���c_����+����p��cY�~達���1�z&�L9g���ԏ^�)�F���.S^:�x����
K��I���G3҇
V�ط�a.��3{�{$�1�0��!�%Ճ~��W|�M��	�(̲���ξ������ei�O���y~�x���� ��FQ��ݢy���bd�]��
7"�&��k�I#܄�`�4k�;6aJVlO/ȓM�Me�����%��"K@���g����������<H��c����L�{!�`�(i3jݭ�F���p� o��]�7p�J��PW���lҟ�!�`�(i3�����5	��{�OF8F���m¡Z���ֳ×�I�+��!�`�(i3jݭ�F�������a�d�tu���ād�,������(]���+�J��U<o^.K�}�{��$&XT
��"{p�������n[���/b��{�P}�зq8�Ј)w�<�_N`E�cvR+��}Dq�f��.��Ԕ�9�JzM�E����F���8�TP��@E�`�8���&�Q�$_���9�JzM"�,�>E��4];ˍH����TI��Ԫ,щ�"�J����2�q�ۢ�)�ak�m6x�]�V���t�����[F�a�+֚S��~��������c����L�{7�ܥ��2�`e7��9��×�>�����>[Hs�?����H�Ud���7,ԯ���gn��Ab�%^��}Dq�f���<E�f�y�-
9dZ�ד���b����8�TPO������=��Z��( �s�٩���I������.V��:�7�ܥ��2�`e7��9���I^Ɍ�ȓM�Me���?I�g{��@���g����������<H���B�r��!�`�(i3�����5	��{�OF8F���m¡h�q��d��ZuH�!�`�(i3�����5	��{�OF8F���m¡Z���ֳ��m�,�0��!�`�(i3�����5	��{�OF8��'�PD��I(��<�,9��8��A�B�r�ݲ��+�J��U<o^.K�}�d	c�b��8���&�'�al��p���}���i!�`�(i3=]A��O�T=�4e=��-"w߻Y��}Dq�f��.��Ԕ^�|n�M�!�`�(i3���D	��U�l>o��|��P�^/�h���/�d����������622���k˗S�d�"�,�>E��4];ˍH����TI��Ԫ,щ�"�I(��<�,2�q�ۢ�,�Xʚ@h���+�J��U<o^.K�}/��<Ӭ��|#HK��I�7F����x��B5�!�`�(i37�ܥ��2���kܪ���*�LNm�`
 ֢����e���W�\�h��&2��>/' kx�]�V���M�K�=g�H{g�q���I(�c�M��r �6,�Xʚ@h"�,�>E��4];ˍH��\B�����g�q~[{Q�����#�(y"BT�(���B�r���E����F���8�TP��@E�`�8���&�r��SQQ���bK�&�B�r��=]A��O�T=�4e=��-Y�VN�=��Zt%��m&<Z�#�j��A������!�`�(i3x�]�V���t�����[F�a�+֚S��~���������B�r��зq8�Ј)w�<�_N`E�cvR+��}Dq�f�]|If">����A���I!�`�(i3,ԯ���gn��Ab�%^��}Dq�f���<E�f�y�-
9dZ�
I�Vd���D	��U�l>o��|��`��	4��=����t��cg3/F�~f��
I�Vd��7�ܥ��2�`e7��9���I^Ɍ�uO	Q�� )wS��U���z�x"å!�`�(i3x�]�V��:�R3Q|�I3ܱ%�1�B���h�{�p�E��.�^,W����L�z��̾_4k&}ǝ^3!�`�(i3!�`�(i37�ܥ��2��4�7S�ʎ����.N�̇��Q'݀�=�� ��-�є!�`�(i3!�`�(i3!�`�(i3,ԯ���gn�M��sMÜ�}Dq�f� �0��k{.Dt�0�Fc�&v��9�z�ɍ�Qk�>���1=�4e=��-	i�/B�,�����z|�jO��8�|q�̑
�B��+ H!�`�(i3�E����F���8�TP��Vch�8���&�5�R�U%GV�<�nbBI!�`�(i3!�`�(i3���+�J��U<o^.K�}o�C���j�8���&�5�R�U%G��_�ܔQe���b�!�`�(i3���+�J��U<o^.K�}o�C���j�8���&��a�O>*�SО�� �!�`�(i3!�`�(i3�����5	��{�OF8��'�PD��1_�
774\51�]2�t��MJT�!�`�(i3зq8�Ј)w�<�_N �VL�(\t&����Z�_`Ogkl@`��m'��r�Nt[NzigzA=v)�E����F���8�TP�WB[�e�^!���}�w�x�P��_�S�
ut�U� ���_j0��.@.��}Dq�f�?�ᒹ�G�7�ܥ��2���\�:�"�37�˱�5dʯ��V������,hu�%ho����G���r�_������ȍry��	z�� �����ˑ��N��k�I#�\(z:�ĭU�A����N�By3��<Z鎬����a�gN�3c!�`�(i3!�`�(i3!�`�(i3�����C�#�ҒIs{m��M�>�?a��:�1P��#K�SM0.����H�������5	��]�!����58*�!�`�(i3!�`�(i3!�`�(i3�4Y�g�~�r�;`Z!)>t{��U��Y���D��L��</Sn���Ӎ�g�cޢ�{l�f|�t�K��0�!�`�(i3!�`�(i3!�`�(i3�;C@����1���S�Y�섫�So#a�VR^��{ӮY�E��vNd�)i��O�q�̍N�By3��<Z鎬�������(����} "m��^�V]��}1;Z�减l|�*"k���(ӈ��4��S;UA7��I+}��[���q\���2��}���GG^'�-l��{l�f|��rs�i���YN���j[��v2ba(􆿳�xE�zH^�7�{_8�Y���˂lq�㜯}Dq�f�F�d������`��N9�J�LQ��w�6�5�p��~�㲡�S�)37J*uc�A�L'�t�O��y�$��g��U-�e�,���6+�#�ҒIs{g4����/�Gg��q�
i�c�r׽v1a{J�����b3�'���Xw�j�7���N�v�1��n�_����Cҷ��e�ˇ�h����2�[Q	��
�Q�}#�ҒIs{vn�lK�Gg��q��Q�pA����^W��k�va���'��?J�J�D�k�7 �:�BF�!���q�%��Ro�����:,:��F�d����"'l��*גǳ̨����2c�8�4��&Y��V��CE����r�գ���^���r�4��U�U~��tn�+�e��j�3����&Y��V�贅����OD��G͘���j)v������Rn%�bM��pK���|�"u���Mei|�J�8#O)a�7�%��S�ғ���X��4tΘl\	�����:�!�uM�����Ի�弳$��Ϡ���"%?S#�dIǏ˨�g����K���=
��P��bE˧�<vr/��S�s~�k<����-I���z�S�s��T�	J��#�`SN�ʡV�l�Y��j3���	� �i/�]�!��5��E0����|e"�@����M��{l�f|��:2QYeƈw�`v@C-�<�6�Q=�Ʈ+ˀa�1P��#K��uṔN��ǋҠ7�	�ߥ�H�^ /m�6���<�6�Q=� 䉇o�M���w0�!�`�(i3!�`�(i3	g u�XI��ׅk��+ņ\.���(b��i��T�ȓM�Me����l��1��E��΍�!�`�(i3!�`�(i3�Q-sH|��������OW��F!��߸�Z�C���!��5�Ǐ˨�g��n&����_�o��C!T*p�VU��Jp��T�����hy�� g�W<��z��}�<ͧ�:|zG�_h��� л��������W!u���-����UY֭���F�eO�V2y/��S:�cN���dt�{�Y�Mei|��Ja#���a�7�%��S�ғ���X��4tΘ���VCS�!-�+_`�������"�g�#-�5�����77AƐ^�8�tn�+�e��j�3����&Y��V�贅���Ǯ0��]㯟B./�<ĩku��j�,�J�2�|bQ��� Ǐ˨�g��F�d������U�We��ǳ̨����2c�8�4��&Y��V�%����B\bE����Kl3��+�I,�S���R��z%8;����v{:��h�k-J����:M���FM�`;$�l���1��in���� zԻ�弳$_N� ����_^%zl��P�;���������t-5S�)37J*u�,�JL���ƍ2���lĊX�6i��{l�f|��:2QYeƈ�	����Zt%��m&<;p�����I�K��d�S�)37J*u�,�JL���ƍ2���l�J�a3mPyS|�P�D�o��C!T*p�VU��Jm�QA�Q* Q'݀�=��&�v�x�o��C!T*Y�{'%s43u�R��]|If">���%�o)��^�V]��}��ł�!r�dN�<@Iv�,.9������:5A��p��1���z\�=d�#Q�
_�J�g�J�LQ��w֚S��~G�݈,��S�)37J*uc�A�L'�G X�T�ys�?����H�c�B���)�g��U-�ee�@Rv����my$�N��;� ��b�� л�d�q=N$,����hQ���}VA�ڦ�c4�RP�m��q��ˑ��N��k�I#�\(z:�ĭ3S��n��@IE�U����S8�=	���/lg������T�\ �́��Wl� -��J�x"GeY𶣂���S.��TD���rs�i���YN���j[��v2ba(􆿳����r
��qő��{r��  <�!�d�<8�c{}�x���� ��6%j_�z��D�-p��n�a���2��v��z�NFX�5�B�ʏ��Z��N�~+�|~Q�d=/� gWVbT+踫g(�r� k�|6�8�Eo(d�J��:��������C�G����]'\gWg��	�Z�kfc&�2����{y����i�q,?5qW�7Q�ǭ�7�I0I/Rxjzӝ���I(͂��-����!�`�(i3�.W��E�g�������(ӈ���m�r����Ra])n#���^a�nu4Bޗ��jw�	���ݚ�Н��
�t��T&���LQ�/81tSjv�!�`�(i3DN��5\����t��PЌt���ߗ�ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 ��׹�3��܌o�q��_N��.�g3Z�7�4��~���%���.�g3ZZ�tH�=����q��tj��x�13�KB��:|۝ׯ�oȺf���1�H���?�d���&��ꢤ�Og�:#��XB8	��K��>w�R���yG�e��bo ��R٠ș����q8h�G[�� 4&Ƒ:2�c<�^<�H+�|����n6�i��<&� �I��s{")8�*If��4�qnw�R���y���,!��ኆ�SVE����7�ٙ���O�Q���*��P�Vr���J��:�����`�x���$y��DcQp�3Y#�踫g(�r� k�|6�8�Eo(d�F�!��c܆�_�[x���F�,�֏��9�GͿK��n	l��Q;�im��ȍry��	gC��� qI�`���-�����1�,��pϓpy%�[T��k��E��\2��T 2����?�/��\��u�7��ĺ�2�a�pn�d�D&R$/����ݚ�Н�����e23؟��Tφ8�$�|�C�(�mWƒ!�`�(i3D�c=p�^&�c��J"O�ڞ?�ǣ©��WT�/@���-�L��Ғ�ۍ�<��W{0`�ǣ©��WT�/@���@hG��կ5����<�ξ�\zǣ©���i�ۑ qL�K�Ѱ�-���ԌY&�xL���2�Y�n!�`�(i3�zsO%!E���tR�/p.0��I�![�Do�9�ݚ�Н�:��+�������4�tX&|a�#�I7��-5��5Z���D:���*=����!�`�(i3B�O�%J(V�K=�u��!�`�(i3�ҀL���G�_�������� "5�]!�`�(i3�M���r��X;p`�l.�	�C�!�`�(i3�'�al��p �8B�@`6Y�{'%s��1ƵS�D�<`�
A�$�1Y�f�?ǉ�=,�ttT���-���*��b=�!�`�(i3n&����_�a�/!O�f�?ǉ�=q�\E��0��A��)}��{_8�Y���˂lq��f�?ǉ�=��ë���6-���+?B�OA��At�&�2����؍��R��I��)���W�w��fD|��זw�R���yxP"�up��%A���h�Mgw�� 
~�F�,���XF:��GZ>.�0����ڀS��d���!i秭�B��@8GS��`˳j[��F�r�f�t5x|���MM
��,=?�d���&�(�6k�4d�kQ�:\��#ɱ��5?�&P-�_.��45�I�{�P�՜���,�ǰ�������Z���zh�����,�ǰu!�OO��
}Z8/��RU��H��<�C�Ar��� ��иܖ��A�.u�r;��|B
y�3~;�>g��4� �㎿���o��A�q�m�,�5�%]����8�B���ow_;O
�J��:����{k�h�+*J�X�$��+�nj�a�0r�uzZa�U2X��������,�ǰ�������� 7�G�Yw�R���yWp�K#J��d�֘u�>݈��Kyr ��6�w5����B�}�R X$L��~ џDq�]ETk/�0��nz�������b�G��Su����*U�:ʽ�fq8*|��@�)s&� ��e���]�!��	Ǹ�y85��3}�@�7 K	����n��,o:%{�7��4<��z��}拋ġC������Eu ]����b3�'���XwKE'q=�D@� ��<��z��}�0z�cUL��Jv(K�V��c�4��s���o��x�8���/�KE'q=�D�]C�:���<��z��}�0z�cUL��Jv(K�V��c�4��sˈ����8���/�:q���0�"��!��� ��]�!��]/~K�#B���7{�ҋX������S8��y�)xʔ���V�� ���`y�����G���Ld�-P�Z:����"� X$L��~T	6:��=�0@���&��c1��v�u�`'s^��>\:��9Km?s�_{X4t<� ).�xg�"z�JmD`�|��K�z8<
����h�d	c�b���q�Y�
p�-�L��m+)q����h��@:S"���E��#�x�&��'�|�7����s�ݺᣄ2m>y�H��{Ф�E8<
����h�d	c�b�IϷ�����q��3[�W�W��<��W{0`�TD��nE����X1'1[��o����󖈣�0F���E����4���N���m��;���g���70��4q(�ٓX�lz\�Q��v�r��Rϻt<� ).�x3l��ڽ��lz\�Q��?s�_{X4x�]�V�����TI���U�����Hlz\�Q��*�N�to6�k""��{��7�ܥ��2�-_��Y�?t���X��Q)�_v����4�F����>���=���a��z>�n�S�� ��,���1��؅��FJ��u6Mn+J����/3d`�|X ����p�IÙ=�H�~�5���l���tL:�C�RH�YGD@�F��qW��Ґ�Yj�|c������l���tL:�;��K:SGD@�F��q`E�cvR+s̮�s�a:�$�77�}�(C#ƀ��=���a��JLm|�Ij]�������K�� ���i7�ܥ��2�/��:M/�V���k�=��`
^8�J#w��(۷����4];ˍH�O������=򩦞iQ]e���}��+�'��r��Zw|�pMGD@�F��qX�ʟ��{ŌX��V�t(]�XS����ڸ��P����؅��FJ��qW8+���+�8�lc��x{�:AO����k�*���t�]P؅��FJ��o�C���j�c��j?;��~X��1J�j�k�;V!%�B�#Kg�je���Yt	�����\�����!�`�(i3"�,�>E��4];ˍH��\�Mb�mOU��e�Ի�!�`�(i3�d=}b�TY���t�!�`�(i3!�`�(i3%Ah�%4
>��XP�����t\��X�i�ۑ qL�K�Ѱ�!�`�(i3!�`�(i3!�`�(i3JHn��z��r9�3���Fz�Y�b>bb�v��UP�!�`�(i3!�`�(i3�Q�^�y�zL͊�q�����7�f�2Y��kک��d��G�P�x�!�`�(i3!�`�(i3���D	��U�l>o��|���JLm|�ׇӭ��v�Ys�S�)/^;؊���:�6ӰR���&v(𨾤 ���8�TP��k���h�%�F�F=��)E]ׇӭ��:��+���f�.`�G����4�t!�`�(i3�E����F�'n�^0o!�[%9\U
!�`�(i3���4��Xה� �f�!�`�(i3!�`�(i3%Ah�%4
>��XP���p�1�q1��]Mt0�