��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����⽸���D��6T�8�{N�/i�kf�!�6��̋"X��:�����\N(h�-����}!���1�����4�0���S��k��Xd�d���{�8�%���AHǚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>,M�Kߤ�A�O�c9b��2���j�:��HA��?�\/��q�k��#W_�0����J杦�&���£mj��̟鬶�Pf�s5��q�Җh.�k�/��HJGS!]$�y�}�t+��`I{*���:��Ʊ�/���"�F|�n4�����zb�-�xz����W�uX[��Х�U?L��}*uT���0��܅�Ü�a�]�Z�!R�OT���{z�n��'�"�>W��6_�I�:�}X`ϻ�ϸ�k���A�A���Br�[����Z!	�D)�<[�杪�9J�98�U@�;M����ڑ����%���nʕ��,�gFv��t?��[2�0%Y&֠b'%ݴ��T8�p�-�g��K�NbM2��_���U����fEe�֩�@��� �B�7��2��X�qV��\M����Qd��}�k@t��lv��Q*�[�3�,�ۇ�v �=ֺ����+l���><�X�e��t��\$�
<��kDD�W�*λy�u��M����v�"&�f��U�'�� ���t俋68|«m@�֯VY�/20�k�G���-�o`u��#Jb6�k`�n7\���n�fļ��IǊ^���)�c��+��=�m�.^���;��?��f�ż�dkS��8W����M^^ZcVǧj���7KT�S� �|?x��8����	��!���ut��w�������m�� �&��>��ܵPE��:�f��/a�&�1�$?i�+\!� lՈ1�<��+�T~��".Q=E:�O��*<��ϸL �����X�����!T Tg��Ӹ{}�H|���x���Â�ڳc�إ�&�_���1A��\��$���  �n�������H�_�	z�&���UM&m�;�*���
h�E[7A̋m`uxiHZs���i��f+,���WF��`	�]=��&��O< U!)�5�7�Ģ�j��/�Kl[xyJ	Vz��F�Hfqz�$ C������*83�BRA��SC���!�ޓ��d��0K릘��vɲ�ܾ`pO�Բp��NV������ ��l�d.���k'�1��O���ɠKy�Y#Ų�69?�~�&T�܎U}��%�^1D��>3<�%AA'u&`��02?6bW���xɨ22�E�+�FUu
ЮΨ���X�w�� \��M�&�Ĉ���Y�D�4�����Ap�l�W�{��f��~R�EbB}�mpDϪ�4����F.p�$�o�x�,ϔ�.~����!~5E�gbS�$��7��y�|�~�L�E׾�zǢ�}ϒY�s�\v��<��~�%���*�/���ǨS��B�����KXX�ۭ����Q0��Ƣ[;��7���i�d't��{M��
�P��Ğ��9��ș)�D������@���`s ��ܘU�	�}5���;q��ez���d�B"�%�Z��0?���$����S�;?,�h��0��B~�<'H��q��D*TP)U?�VzF��� �g�|4ƞ=�тN��o$�B;?%@��K�J؜��V$�%eܞ>5Âa���ie�l�|�G��Km�Y멲�g#�#{-Ϥ�/���dk�F�b��wp6Ȱ�������\�j�?.j=�؅-�K[Z�K�]˂x*�[xIұ��=o�\��q�#�n����E����r��v��gM�!}�� �qysνo�L:v��؍��+,h�	�4�=�OKi�~*�_�tȰ��~B�d��o(b��^u.�'��U�?���ПQ��<I�8R*�Vdn�/���֔?�"�!�����lm����W���"�?��=�[6<��ȅ�xR���ύ]��s_����.����C�,�ښ�n��@�7�8�};���r\l�Go��n#�E.�۠~��� ̣��1��}��ߠ�������+5���\P�U�����e�\���T)��C�ӡ���
���-d|8��_��XZ�Nb��iu����8<|m#���� l�E�4Kb�9���n�>�9$-�0;��gO��LV�w�h0��0ʦ��Ů^��^��Uy�4x�gz�:� ��ʘ��sAĶ.�:��|!y$AՁ\$Յ6�В�5[�_)��"�e|���&��uj��L����Rϩ��he���*n�!�H�(Ҍ �$��=�JXfH<�C��p��.*DtPc�7�w޶B�������\��If��+���Uכ>��W����1���s���n�]��ů3�mj��8���L���ʊ��m�1�j0~��f�m#�-y��t�;Fd�����Y�YKq���	�L&��E7Х��f��q"WhI���]�\�Yn��34�Q|�ݖ��uzs�&~��Rz�g�˔+4�����'��%�u>_�t@Kl�X.���'�_,�JNmy`ʑ�e��*�5�QU��Z�D9�-��Ve�[G�ႳMǮ:\�s�)!ƾ��;���n����hJVU���c�Ѭ�Д��K`��np-W�?���6���x�/_��g��E}�r�\8��šC��vp��j$�Sd��Ӛ�?|(y+����U8�sH�������Kfh`b�)����cY�P�R�{+V縉7_���T\I7R}�+Z^4窫�C�ul�
��?�S�>@�^.��=�},牘Hk���E��������V���s��c�N����>T�ts=h+�sE;��yY����):�x�:������R����@5@�@m�-�����ʦKX��]b6�{eHwm2>|E��\'��Tk�����z� f�|_p��  ��;JvS��!}�ٟ����wCv��/�SWj�f&�l��3�䥁q���*@�"���W:�fJQFE��L�j"����;��c�q,};gq�8w�C�騵���zB3U��6�պ�Q�P��_�{��q��XԬ
N��3U���j9����d�(�_�؜u�`?0t�<k���V$��(��,2�\�c\��7�p���03[���D����ؑ����g�`�r�%�`⽦�|XFcQ��sS��,T*���clqߦQ`�����![,�������Ч��.�%D]��F���RV7��C$A�1#߶�|��௏�ۄ��m瓷��"�|�]s�*Ǿ�s=��d��(!�Ɏ�	����~σ{�� �a�pV~�)�+c��G 	�bQF�޵GO~S7�}��٭�Es��F:�草�|�13��߲0�i��n_�C	H�*����ۗ��8`�l���O�F;9����TC�K��&�{'�������褭����j--��m��\�pd/u��n��(L��^A�����g)�e�Q�6�gZ����9&�X�KWY�s�ҝ�l*}�4*u;����A�oj��kaл�x0q����<)^/����]4f0����㑐[Z䙐@�ީ@3a#��� z�DW�!!Ŝ�ǐ�G�	9D�f��$�|M�4
���w-�}Z������ٯ�uE=ߴ��N8��L�9�a5��oXc��%{,�ٓK�Ǡ+�>�麩5vk w�#��B�����-�]l2_��i!O��^�7�����~l�jo]�j�Xl! ��=�D	b��k��[
���b�Ro�-[՛�5�"ߚ�Ri=�9gT03��t,��cۛ�ց��O�|#�� j�����w��r�w�XTR�٨Ӄ}��n�r��mm_��$�άⳌ�iP-m�������8����&��g�A�T���6*{�L���(�8X�#����Ǽ����T��GO3=�ts${���N��ü��ge��V��{��q�_���3?��t����ء��.x `nY�#k̲�:���u��J�$����s�?E�����ۨ�"�j=��K�؞BA�6��)"��o����6"��Ә�y{��Z�|� Ï1ujb�K�����z�mo�e���"�.6x!��a3�w-�sI�ǿxX��*����뤶�k��>*F"��L������Q�t}��9!��0�}���p�Z�<J͟Ϯ���N<>�ª���u�;M�^@���YS;�գ��Q���1��J��VD�m�����O��('� ���L)v^�4�����.7f�K-R \��N
�����0����)ߪ#$�i���Zb]>��C�-?�X]n�_�M�u�J~\��ec}�MAGK�3��*�I�2�谾��������r�vǿHh_���C�c��Y�#d�T�V/�>�(��43V���;N�����$�Ke�c��JVj�Ǆ2�eL.�3/?��(�n�~�ھ��(�?q��;,�+�	�m�xS��H���|1/����"i0a>��/���X+�h}�As1��N(v�t
?*x��gBB�ϻ{�i�?���ݽ	�r��΃�<���6=�F��1�S�!_'l�F���� �����d�Rf�����ơM]��@�/�π�%�!6K�?{��hRd̎" _$_�W����-��Pߧ�.G[���?o��?mb?"L��)�L���7���1i�B��W}�k�� þ�ZFy>G�P���e.[@�`�Z�:���-��3E��E��g�͈UXJ�������5�CQ��V� �Q��4k�/�6�a�@��t�Sv9EE!�Uã[����x�f�H��A���r�|{�;�ƥ�$	p��roD}���:�aT�I.����|�G�7C�wd��ԅf��K��~P�n�e��p,8�F�0X�Zf>��ԓgӱc?eg%�ߛ�2S�2i����?ɫ�)��ky��lF�����nruvaHL{bb^^�W�yt�g����dM��>~��$>�E*#�7`S��$1��.Nƫ��f�$Û#��Y�j)��^� ���i|���&(��t��B��5&E,au�aI�\xd����|ndM	b�HOc.��`�/k�E2\%�0&ghKk�,���Ӱ&kq�T����II�M�M�&�X~ʆ{�(=��ğ����UV̌Kz�@;���I�k(�H������:�9i�	�)u"�Ζ��j	5r��Ӕ<��L�˹�CR�06���P/�,G-6�p��l�1o�L}��&j�۹�W{�ۑ�#�����?����lCY���>1ܢ*��󘒪�Y�~�>d�У$��2V19w_zKlt~R��_�x!���a�����/#�������t�s���D��|pf�ؗh��V�!�#����a��#�N�����"D��'�T?�B����C�&�#���VƚFǂ�
Gۊ�Χ�5�;�����q����p�M�t��Z�x�p]�$�w�:����E�vD���P���+�s<}G#��[Q2�!�\�@�fc8��W�%{ܛ�0���9X���t���-�ɨ�;��������m�7}����NV�<�����l9~;��Q�c��|��t�����T��5��L-�3���+mfd�c����l��W��$~Q@�v���@�A7p�+�R%��u?u�)(���>(:�=�Ҧ�Hp2��&����I��E_0h�Zӓ׸zA��|?{G�����%�a���S��'���a9�rw�U���p�{ɫ�97�1ϸW��g�*��d�!���P^݉RW,Jk��N-�Q�� ���G>ƍ4���4�UuF�?��=G t`5�y��c�r�|�Ͳd�����u|S����Bb�tvy�D�r�+���iLإX9ϭ?I��5���Z�B6��c�CL�A�G0m=��;�M����W�o��bN��4n~��ڥ�G΢�2����\M!鴴�9�����R�E��=F�o�G�PZ�
��*��A��	(�E�>�l��Kp�R��Lx�օ���x?wK @�P��>���Tvԇi�F��;��ju*�:8b��jkg�;���S?��ї���cqv]���s��m�Ir���W���\������W��ܚk����ԿR���
Gg
��-x�?N�����ʚXF��dB�b�n%l���a�>W�{񵍎O^O$\��am��K8����pXTC�D;U��d�P
���.�4�Tl�h����	�F+��I�I�B�:����f�É��ZvB�c�����
�~�T��"���/m��&����Om������r� ����e�e!e�%_�p\�N���-��o���j/� ɴ7U�d�����|�0ew�g1�]v�؉�������ץ�2�+���v{G�ߴ=Gft�'�z<Tw���-����E��m�ظd}�T��i6��r�ǃn-O����M37�K%�f��s�-�{��������]8W�!�j��(�n��p����a:�:cdj>PDT� ������9�*ڼΈ_`_�6mC�\A8�B�Ԓ��;����Ic��T�� 4���_hQ �(b�I�;�g_P��N�h�^=�sN�c��>��}�$�nH�]w �������bTx.�����%�u|�3�BsFC�?�?,O��M�2�Q���z���P�ZG]��G����dP��q�t�e�� �a@
��ƞ��4r��zi����kg����Jk�Ŵe�|��,֯��w&�oŁ햔�tVw� m�c6 K��U�pr�M�� s��˵kþ&�*W���j�x�6s���x���	uv�O�|�;Du��i,��>Ni�������{j� W��L�aa��t������ɲp�T׃?�85�[L�)�-�=��8ta��o���јy$tT���8�}?R�W柙s$���]c�	�\%�]�u5+��č����[ή��Ӫ������x ��w�[Y���LƼ�?�%!7ɸ�\H��2����nyl����l��vq��k��s=L�͚�����G�
蕛�6��5�'&dZ�>Ɲr��P�[���B� �TH	�W��SB�ˎ5�P��j�2y�/���u̬7H&cW�ū��z�D��ɂ�E�Y�Ѱ�+B�����J$�L� _��>�cN�[��{_'���袁N0qe�����)�O�M%��!�����P��΋!���� �C N,�yGc��Ϲp����v���P�-�H����V��Y�;�G�BɆ��e+��#a�%@7�ȯ�L�!�f����N�V	gU��H���qa/(�@��"�2O����x�(��C�4�����{�g�b@��L�p�c�`�K�D�����ƣ�H�)P��5y`v�݉/�i�L�Y҇�1�ݳz�D��*���ײ��z-Eɽe<�P=�H�D����*�ȖU��h�Z3֝�h
a�2#h��倳Š#ֈc�lZdvB������`)��6I���Ĩ�J�����E%���8S�����y�k�f]ޭ�G� J�y��Ig��~��'�X�`����NV�(��˿��	�|�ϡ(`Ŏ�#ؑ����;BFU�vz�q&4�]���%�������i~ˎZ��Wa��Δ��ޡخ����[%z��\�p�����Hz�>ST��#�u��sp�w1G�`�=Z9 Sv�]2��",��+'���\����D2ri<x�Z���'��c݅�N�=�j���Q�O�s��Qf��z5J��ܐ�KV�*=�����Y �����g`��a��:�
���xb�<����jˋ�(�fQH�G��s�<xhwP�4���8�d,i*�swDK(@�C>�o������< *�p[<f��L���ir	i����,�/p�R<�%<7�U��l���j�̍7���듂�J��l+���z�IW0�3h��ҙŜ�����ѥ&��h'�>p���T=>�����ޅ�1u�~ϓ�k/����!p�ޞ>N˼�2wڪ����C�D����O��G�E�ѧ�e�F��oj'��� ��,#m+�3�공��֠�p8���iC�%j,�i�<�e������nٛ�[��cˤ���)��0%U�\>e3��@iq�‷uߖ=��� �b�\��1��kl~(o�^��l ��y��__ܴ��e���W�Һ�ҕp�ۉ�t�kX ���v�uh`����u��D)��%S��M�</t���6&��pu�i�?�>���+1Z�wn����4��Ǜ%I)��A|TUk	�կ��%�����E�b�>�h�4��a��� �"����{�6x�UM��:����S��u������|�{ljOug���k�!�ϣ�ɶC��Z��b�,�|�$��t�{3�Mg��k�$����3!�(�$��֌���|����vkK�#�ȉwIr��3�d��C�z�A��T-�iB�p�TRV~��X!�lޥ���< �kE8?�L�1�gV_���0u��+��k��`Mh��aą�R<��C���qÐ�KLw�ȭ�]+�
t7°Q�D=8��w�N�n�墓��[(�
X=ZB�)�.`*zǰ��7����qӋyL5����j�p��1�]kӬ���1.���(P=|_K�f^c�>m��XP��9��B�F��7g� �J'��pA>�QvSOI�Έ[��0���v	≆�U���ʶ%�ͨŞӟ��r��c�U���^�[5=Ͳv�/M� �K�P�(��>����$՘l�O ��Z�	��1��m���n�iL����5�_� ������8��]$!�����ҨXi��tYf�;�Љ��v��$(���BqE1�jk��E�%�V�j��D]��)�D��Z�K���2��z߭�#t��������!��,�Ut�ו��]�}j5�DE����VCc1�����t�5W�g�W�����ehk��"�,n�FJ��T��m��gڍ	a��/��)�a��K�RgE=_M��L×����e!���~Y��ۂ��ЊQ[s�P��l���Y��t��~6�߬ӽ�����e���.|i�Kic�j�_.	��Q��j�M�:�R��u��[�j�[+�w��B��e|@"�Gur�h���HR+����S�� �HM��^������6x�ϗ�*�KN���t���2�2��V�e�/���:j��b[���Q����6;	T�(%M<z�&K�^]'���K?A,�!�h7�!G��S�5��¼�ɕ�i>k��"�y���c]�n�q��3�WH��
��"��(�t,����NI�q��(�qu�DUz�����!Du{-Ի�Y�k�c��cM�:lv�/���3�x�$Ys�Z��/?�d������2����V�F��_�͈��ѭ��A�2�aUK�������C�AX7+��QK�P�1Oz�x�[q�ư���f[i��1sgz�7��N�M[O�Q��;���Td��=O�Q���$�Y����Sp�\�5��?B�hF�?�p�8��=�f�.�x�����#/𕙻�&�"��kU��>��S��$�2cʶE]�p�Ơ?)����uN�"�Ɛ��D��+���4�����<�)6П-W��ԃ�@�\�b/VO}����1�!ٷ4gh7�']~&8�+I�
�t��-�A�C��Q���Wߞ@�
��5�BΞ���seɶ�[V���߫0���^������1ѣ�����F085��H�L43���v��U�4�'i��25��MR��k��:�)cI�`qw�ޣ����>tZC �f��j���?b��W�@�mJ?l�U�6�	
0g&oߊn��ܮT���"��'J�3�k�m���g�[�J۟u�|r^���<H��N���*����2� ��4gCS'ߺ����ē7;D_۟�۳y��u�E煋d�z�ul�oj�X :;G��)nB
k��F�\��˃�^cO;��\x#L7��=>��neCZш��pĤ.[@ιE���P���*)�CqA�}/�H�-�W/�m����6P�(��1W!�_(�mФ;I�h~�Q�(�=Aڔ���ߑ9owdXMZ,�l�7{�1X×u��Sx���Eϊ�d�3��[:�� E����&
t�ޮ�;צ�lnX�%i��+�:~����db�
t��<�XG�=��^�g�0TF�nW�8N@����e�wue##F��������������0��I�	�z�nU������#�����%|�%|�Yf׎H"�"�uG��+P}�)����lGD����{g�Ҭ���W��`�<)e�4]�5 ��ͯ�aծm�^�YֵE�H���p�y�I���v���V�'����fM����b��埅���z&n�Q�ŐG�nΰ� )���<-tħ6
sbD�&ҵ��w4jez^'��Iyke己��CϚ+���۳�Nۆ*4*n8k�cn��{�`2��C��	�>bsD'��lU�#���|	ǁ���;�0���2?+�����`�p#h���������A)$�U��#��Ԙ�}Ml��d�O�ci�t��(/]�<��������K�x��Z� V��\fԔ��$��Y�.�a�#s_�U�QT��j�BR��~��@	��c�%�=q�Z�X��i�%,�^�nocb�@;7�x!���q��Z;��[���0������u��FՌ�W�Z��>_�ys�-�"�.�%��^���d}�RB��E��v����u�XO��K6Ō��VM�k7�&��֕�$�P�Yq�(����׍~�z?�	�C D.g�����9���|����b�'�U�n{wq�z��Q�~�*��}�5;~�4`�y��bЍ�͘7ש��%�)$\)5%��Rw��c�3��G�&y3;�7!=7�0��6Mz����1-Ik��R���\�j�NКzs�V�pw���g\��X���[0�*52�-�;X��^k��ZS���4Iz�<3�Ѳ��'÷@�&�)B���T��<)� �W<bZ'��~���v���	��Hw�(֞�Pi4���e}�/!��'w�x����H�r4GԻ���7���6":��]l���#������(���J�E_
��ǖ��e1�S�	��K��D�r~� �����jބ�{��i �Fǚ'��S�r��Ʉ���	#�9��G�ǳ���[WR�ᗻ1�/GMkb	Qz��2�wN��Ti G�����i��ʋ�!M̽������"/t�kr�7����j�0g/�0�	���
!�&�d7cUܾ!"�a��u�LY�+���T�� ��eQ�EeA�-�O�aN��e;��M�Z�����eb	i�svn,�+lHH�j����GC����U9