��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����⽸���D��6T�8�{N�/i�kf�!�6��̋"X��:�����\N(h�-����}!���1�����4�0���S��k��Xd�d���{�8�%���AHǚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�A���0>�kz��/ �_M��<-�[a�%�����'(�S��jS_�,��8��T�.B߫C|��N�(ݝ_l0fS!��mYԥQ��DF�S;���h/��9mϓo��ޗ���;,=1�7�\ŧ�Кb�X��IM�i�+F֗0UYz�!�K�y]'z��D����;޴�&�y7동+Z�D܁Y��t�AT���Q��<��Ѭ�RBb���Z�_�"u �}��޳`L5�Us�-�����ǿ����x�ze��}g��t�  Z�~l� T`H$��U4ɧj�P��[�?f��fZ�W�1�	(�����zi�q�ߎ��@��}�K��Cm,�\ _�s��eÁ fXg�ķ(�5)�O�ۏ��j�1m��p��N�?,�Wp�6���3��!uD��8�P�y��6A%3;�:7�9��NR�V�� "��4K���p+@���,���}>Gw=��`p}Jr h2Pa��#��O����j_� ��9�M���ˣ���_�S>b�����;��mv���đXw�e��b@�m`�<�ҟ��?=,���Y)r���o-�`8/���k�����$%D�4g<_G���e;cr�'��/�������jC�ȊAuu�����)��b}=�N&<~�KblyH�^��2�u��к���� �#WqP��L��8a��<�q[ b�!�s����>nF�6�.�b�=��ux�{�4��a�"B�/Z��Et0�s.|�K����>�C#�ˑLvC�.}R�:a���3��{�;f�����ML�mo���3�o9�&��h凈��4�T4`�ɩ(���|���	����c��jM[��^N�"JS�1p �V^@�H�3/o]i��H�]�Zǻ'��L���݉	�w��śT��k�kޜT��[#�����L��׺�1��|b������!U��S�T�L?m��t�v�/F?�7����ujk�ADa��l@ƛ��AZ��W�r�j�W�!����ھ���k���\��~7m�y�eI*g����]�	^���/��?�Wψ$��c��|��>\	r��W�5��+ƓҜ��D��a�EZ)VZB1��x����No�:�3;!Pa��%|�t2w��\�����I]���y�T�k����BB���,���cJͽ?��0���`�nJ��t�~��(��ρ�88K�}�Y�e�c�N{�j"�.�{��������`���jb�nfT��침`�|5OR&=���n#��b]|��M��Ot�{,����!�ׅ�	"8Lh�+o�kw�]7���7WR@ �jp�=o�\lj��T�p�Z�?����Kh�k���[�ͷAG��/P*����B���`��<{�-S�@�y݊�D�*7��4n8�aUJA5��m����#�ǂ����Z�~[	� ��,��2h�ne�b��%V�]��i=�k��,��*�|��sl���.��N�_�y^��5߽��bdyy��B�n[��Īq����;��R��i�V\]�W8e�Y�6ew���A]�y/Z�55A�������Y�ػu���{�H�x�{�����s	ʉ�F�u�5е7�rT�����=l����� ���gv��/����������VprT�x�?/�b*�T۽�i��籏�2o������S��~A��0��j]�L:�s��%}�=�-WOJ]��+"6�*K=)����ތP*�/�ם�p��""���T�J��?P�3u\E#kw��m!l��5�`J���.+'�\T�u�~����p��/F}}���o-畱%|���)��u�t镐�=􍫗��A�%�������P�*#m�T�ٽ�qf?�ԟy�:�0A����G#�p4�㗍PoA-_9���OS̄{���m��8b�3ᇽ�If��>B��m(X�����U"�_�̏	�����O�oIB4d���y%����S&O�wh���y������R�o�J�%�';�Nd����v���{���G�Z'��O��I�1%ͬ�C��4����t�㹻�e�<��������=���1s�s��]{�w!z ���1�9�e��Y@0�
��K�i6��@�v) YBY��ӂ:ڐw74�z��+���.��+��s`���y	�t�+A��u�m���I��~��4Ѯ�_k������F0���fr�h�tDQc���;Jm��g#$�'g�{�>Xy�C�6�=�>�u�q��(��.�����uqց vv��G{޳E�Ow�ţ�D�Q���|mN�*I�{b����<%L2���z��ܛ���By	��m{�_q�[��E�Vk�����-�*�X#��}O��:.{84�]즞��<�L�:��Ε[��K�JxC���3��B.N@.x ��}Mvo :���U�ɍ��\��S��%Lg��L����Jh��E��S�����/M�� f�����Mk~�ּi�n���vG�sI\��g����S��^N��q����x�YC�8	}�\b��]��)ৗ�W�̥��ZO���)�����n��{Xf���2�&�A�
=W0��Tw�^� 棸��ϼ�B+Aji��'eG �Yc��P�����Y�� ��_V�wRnxj�/x!���3�辴>�%;K�!�wy�W]�jz��+��vP|
���IK�"e/2G�#�w%�5��HP"@ mh�%�<b5(��d0c��� �vpC?i<�������`Xd��hKW]���������-�d
�!>�w�ת�q�H��A;�@m���v_�'���.����~���� �W�B�_�#	�Ys�=͚��s�Ll?��z��i2�qKߒ�c���~���ו[��2J�6�F���l���͖�u�}�*�kǷ.E����Ȏ�C��*Fs���>�;j�XY-w��[�%�ǟ6�~��Um��/A��S���������4.Bv�Ck������/)w��s8q��;+Xv�B�U�JwR��a�� �_����9�
6Y��KIܖ���~)<'1`ǉ�D1��e��[mG�	%EB���kO
�!!���{!�0��k���&���~�������_�xӎd\2�j4�к<١�z�b68�� Z��lRE1����l�9%L6�b�_1����1�y`Z]��SZΣ���.�o*&nc��e�H��ޚ�pP(���2�hR�3-Σ5�|*��
�-�#�lM���Ĕ�����,�G^1U�R_�O���R�x{U�Xheѻp��[�p��R���6 no�I�d��7��V=�s�޹���09����͘f�=�r1p�)�)�n)=DE3�^(ޔ��a*�^�/� R��,��~V�up����X��>c���'���������hP>�!���m��ޛ�w�HB�D�}�(�8�UiQFu��w���f��`��pb��(�u����D`[�4
={ �(����m��n��L��/Ȣ�Y5q9{r����Ŭ�
Qj!!^l�PRn��m�J$nhQ]��&O������׋n�s�Ɋg����-c�<���[��ca`1ށ
;���!'�t�����aI�z��*�4�t�v��ƈ�0i!�'���YIR^�uh���+�6�qG�m��*:}A|����HS����2�:+�>T�on�1��x�'5�T��An^R�n�_	����Qc#�\\��H�#����?�ޘAt)��%���� �[��@�|�拿�o��d�8�3�{���W����L+���u:ӅA�����tXen(������P�-[�],��;�s�a�#��
��">MnG?���q�e~��8WZ���Y�9zF�Ŷi%Xr�F�%�L��,79�@gS*�[�L��f>~礰��ɍ$���e��~f���	���y\'�C�$C�E�9��9N�e���-��7���贌���5�y����u�]�y�zu����c���M���Z��T�<��!�8�*�h_����V�z&����mc���p��FV�{���O��©�x��(��ӿ|����#�#��L��X=l-��P䌸�dJ�"�R�F��hC��uMNׅaX�Խ�ߢjGl��8QF�t�k.F?b���g|���G�)�\4"�
��x_��YQ3�!�>���)qM:�>^u���ύ�1���
5�Rb�*h)=�Iz�&=UT�g�p`�uh��T�l��)c;��=�Tj��ƌ_y{0,oK��ș����yn�ZQ�RZF���wm���d�0�ᑆ~8-�2��m�M?�T�Մvm��R����Q���2�f%gI�GG��<�Җn�����@�^}�K
�}��+`�6G�Ֆ�n)aB�`�/���(lj�z�h�pH,�{���HA-��?q�u?��q�П���ޟ�;���:���8�E�g �s%���XH�e��V�aU��UFl�,�Mg.3M�b��Q�����8p��%@��ڛ�����{?fF��"`�<��3�~~�o$�ؘ��L�º$��a���GF���u�����FM#l�#�ﱢ0�+EH|���lm�*��Vhn��8~�i��a��-Axd� ��/"5���7r��a�j���>Vf���=���ig=M~�y	Lq]$��Z�w����z���#U"n���I6��澰l�3��`����`��<�,�8pG��Y���C�h
�����w���Q�S���iE!��E�)kw�t�-B8h!1�<��ȜA��w6/�b�'�[&�Y�r���갨ݯ2�&..����J�^����8i�_�!y}��b5J)��.5~Ū��� w���X? jL�����d�F9)�6ǔm��UK38�I)?�����Kԣ׽F0�HzFZ�J�r>ؚ�-Nm>X��U�Q1h��b�i=�>r�,��Na�D�~>�����fQ��Ə�F�P��NݺN� �vE]P��y�+h�m24��|� ��]v���?�Mwr��x|J��Oww��C#�3E���J������F��z<�>=�1�����`��K�9�<J��8x��Ǡ�6����uvc�&��C����}��u������[�����Bfjl�s`��& <]� �^)�^h���Yd`��p0_�|��B3_ZH	̪O�1L��x��0-�^ 3��j��6Pu�M_���,�Q䬁�b�#����h�̬+��������J3�����Y���)s�	�no�qх�˕�W1��~�q������]��*T��f�]OA��j�?x؍��S1�~��@W���qf�"�X���K�ַ�C�C�"����g�lP�$��>N>R\�u�n�;�Dm��nG�x�)�]��(x|�q�o�$ϖ0X�?�MD�౹�mp�cCj��z�0���QV@I�l8{�j�k��k��a�o�Zw�:a��^g1�eX�`�tN~��-�C��j;6j�����JM'�����l�]�
1�%��R�yj����X�y�[�a$�m��e�`�-��3�H|smAx1�쟂�8�H�(�n�a�K��6�P Zn*&���WL^�7�ͅj�hX��+�ٲ��x��y2�0K ����8|g�mb:�@��9��e��n�Ş��'�Oj0c��U��}i��b"Po�b�Ha9�A��UH˸�}@7��>�����W`Bt��'ux��m���&i������⧷�T�^V�f�O�9���8���s���QW�¨l0�]_��$)h�lf�������[�3d��.�@�W�I���A�� %;}n.�t�i��5��
H/)٥�"R�����C�j����B��x�<4�+i h�8[�{u�}�
���Fs�3��Ѵ=~F&4��+ې��ff�xV{kɊ��	�W[����62z������
a�����ϋT"_ t��*d�=���} ��:���,R�Lew�hc�Y����d�F_yo�e]�'!-:�\�;��[��?�S��2���n�Ӥ�$�nX��b�o$�a�Ox�:���-�_���4��(�rբ,��0}	kBU;6j&2��s�iP��@o����&+*L���U����e"WY%6��?�(��g9�c������e,��lD`W<����.�=A��2%�Ԧ'�,=z������Q"OՍN��C� $ai���[z/Z���Z���Qr��,I0� wwq^qܞk�{�x��{���%k{�|��qO[�rrsu�%j�Y�&�b����ݰ�KΎ�y��nu� ���s
��>�<�d�yJ1��I!�ȑ�i�����JoPz�5��k��(<?U'}^���q��W������ɯ���4�������z^����'����@�Ne�� ��n4\\�Oͬ^)�*oit&`h��
����:7$���͌و�af�$ׁ��Y�A���Qh��O�D�+��x����M�������u�CH�Z+f��)E��pw6�tv��;]�^���A9��l�	��ܔ%U8�+��mi�����#*Ӑi�>a��kr^�!�i*�����R�y{�zܘ'E�<i���H��n&�	j� �u��ǐ_���բ =�֊h�I��?��#����~��~rO���`����#j^�x�k2��ȪB�l��L�����(PC����K�x���O_�^P�/3Z>'���aZ��u���r�f�������#�x����z޿�Ο%Jz�Sj�e�Q�,�%�F��A��L}����m7� �^<�%Jg��UO�_��4�J�$k�&�e�;*��7�h`MMQ%x�ha�V��5�u2.�.�˩�X���
������ݽыc�,��;�Π�m *؇Y7�({�c��|%���%�5[���>c�O�n��ʶ���0�dA�N��?]�%�v-���OS���I�gcC�o�S�_Qfzg�#ĭ����6 R�����1��\�"�����u� ��	�C}���wG��`v��f��+X�Bl%�ڋ��h�*`$Q�:)cm8i ��H��ZMu�!`�B�COH����H�#̀K���n�"�A�/��Y�
I�Ç�>5������`;��"ϐ�7����(V���1;ދM�-=(�l�1��stp��50W�=���LJl�`�#��/ۙw�t�x���4Hd����W�J7'���-F��'�_�W��'������h�z����	ō�r�:�]���w�n��n��!�)����w�>F��Qj��8����������*b���A�%�>׌5^����^����S���>R��٫�����,cѽ�~g&�ҙ�@iޜ�iF�\-�+2:��-���;���*c="l�mV9�7�4�о���>�W��䵎���2r4'=z�)���ӊ\���`s��B5�����^����neIE�St����۰n�~���������l��)�f�'��@��Bt�Pxi��̳�?5q���N9���؂0k�P'ŏ�.��n�'�Xp^r�YS!���������	��r�j�N�h�rcCѢf	��gr
����/AE�'�V�u&hʁ뀌�Q�?��mT���P�׎��Q�>-w��(~J�ܭ|��ג6�k�&�~wM)r���e`}�+�%$j���ԉ���ȏe��+N��qd29t׿�H�au�Ff�;��S�I�qٱRV�<1E-�$>����2q.���"p��U ���u�r�Č�q p]�$�O���@0DՎ1�� �B���:���bp}mo�ѯ}�3�[{��E�Ȧ~�zT�$�ѐ����8lwΥՑ��a��)9��h��Y�^�l���u��ٯ����H��x�J
�|�h����9�T����Q:�R���]��-E��\\Q�l��4Ɇ}��"�a2�a��K���xa%�� ?�q�|��*;9�)f�I�(������H�eÆ�G�/�&�����7}�z���2�r^����i��?LD��4g�7�ʨ��W�W�m��	9_ bt�4�����ׄ|+��[��;N�\���*w�Q��h�%96��ȬTc�B:j���� ��=�I��Ml'���ӭ�ڢ|�%�j�  ��L䘕��O��O�X��)��H�8�h˅]��}C�w&d�+�C^	�������c���@f����O��3@,��M~�<�X��N�c��X����K[�.�#܃���ಓ7Ʃ�Wz����f�n��|�!&Z�m�-no����E�ڃ��Y���@{D ����qh��'���ڔ�W )ش��p�<p�4>=%%���S�'G�eע��"�o�,��:�OoM�0t,y?����{��S5��k�����$������V�)�e�:��+v��!���V�:����ֶ�g8��{�j��4c1x�s%k������;�l4|=���ڏݕqC)�o;Yo� ��{X� wOU�б�x��^a���,�s��ҩ��`�e�+�*p�`U����Y�u�|��P�+_q�L*J�n�c��,�GWP�/�j�H&X�x��Q��(�)�@���__$�Gy��?�Ȼa�g*C���ݮ���N<9��y~�~4���r1.�%`,�#�sW�o��L$/�6!|Ae�&o_��Tĭ�Q������w�ۯ�����<V�,���|��l�Z���)p�kmB���ւ�U�@�ſW��/*�:kuȢ��ǃ������q�_maVJ�=�&;yq_�z�Cs�;p�B��	�>�_G�A��'��=ꦏ^�Y_X�R�H�^��sx�K�l����*ƺ1����ڦA`�t� _�
�ޟ!>��5���8��@`Ha��C^H�O���oԬ}��\�A�d�{�B����2'u/�ƺ7��K�Ib��m��i{:2�{Cs���ӡ�A��)�`�oa�ࠟ��;y,������ۼ��uL���[��;¤�[�	�02
��.qJ\az��1H wfU��"�F:x�hO�,�~X�I�EI��Y���2�L�>ٽ7?�L����f�%+p[c�Z���YkR1۩[f�5'��χK�{ˡ����S�kߌ��.�vH0M��MH2�LG���m^E1���}��b\"D�J���b>`"gW�������1�'`��םGD�1 �\y?�;��j�#�mC�Y��B�?��P�A_z�	A���݆�h�sU�='�׶��
4w���C�Tu�f���}H}B8���4BuGZ�.�c�{�38�ƍ�3�̿��ͱٕE���j �?�#��㴰�ܬ�� �#tz�f���q���Bŀ��5�r���b$�IG�c0�6� ��r��<_���V����n<J��>tqNTp��{6��@E���(�M~$�o,ӧ���N���K�vp/��AOĆ���>��W~8���9���I��س������R@���D�QbH9t:eU�p�M��Vx��u2L�}�`q��]�=����"��w�r;��x�s���,�t��Dk�V�G��ru�<�m�:QI��7��80.��A }�n OC�B�ٸ����X�rx�S������Z�ꡮ���y�Xn_�ġX}3l�'^ɇ� ������[�����A7G�����H�Y}�K��Ć��ւ���o]a���sZR���^����}m��z4,	V]��uLz�M%�{n�>�:W`P�D��Ы�c!#+r�4����' %_�č)$����`�Ia��r��zX��q�Q��Y�:��3�LS���]��,�����z�'h�<H�_�]_�#��/�?!�-���g{qo &����>)�����������2�@Q��dwԖ�k�+�7�{?�_���ܚpfzMʝ�'�bC%	�<���Z(�(Ip��4Z��S��"2h1��N���[�ͮP<�z�	^�)���U��
�u&���qS�_�fE���
8���3���Qt[��o��8�Sp =`��9�<�zx�-��J״�d,C�ڧ�B�yF�,��b�Ј��b�*�W��o^� ж۳���un�^�
2 &�N�az���SfTy����A�f^{�=���i)7�ު/�B�|d��B>Zt�kB��O�
b^�p|=T��ږMcK��L^�P	*���"����a����?����y�y��Ҟ�d�3Ewi}F:��Ga�����,c�V�S�]�����B�ϖVQz�9/8�?R00h���L}�h�k��4F+5�F�����G�yAa����Ss���FC�궖�`q2�Q:�[t���~�SxD3��S�p��Y����
�9+�d�'�J���/B�l� � 벁�#^��FZ�v��%}��I�^v�ґ�&��
9��M*[ɻ���|�+�+V��N�b�8���[O���%�߼�;�J�Ỹ���~.�,Z�+V���C�=�� ���AEJt�_5��_#�����oq��·����=��y�|��{��`񧪆������>1M���U�7�l��E�9a(����??���}�5���	sa=�����!���GLB��k�;s�aI���HC��8W�����O˥�b��y�#�����u;11&!���/���b��!�*^��ϠAN�4�ʯa!�H)���'�H��P���M�������%d<�:dB>��~����>%p�y`)H�r����D �[*0�5�E�3.�'MV�	Ǿ5��8��(:��nI�Y�9�ba
_��Q�*B=X�S!�^�$Ũ(C{��o��L[kY�B�uV�̵��\Q��-I�2���-��3��@k��%���ŀ�b�;�s!6S��9����V�;T���J�AM��SC���|ݠƟ;�9w��S�NL��+ 3ԣ���� 'i���Xsk���}O���^k�Δ��& �S$�nΰ�M���ȥ0���}��8�� 5�^�]��h���)� DS�T �ȷ���*���9/)�^"w
�G�����N�T�H�����D��9&N��哠͟�v��S�