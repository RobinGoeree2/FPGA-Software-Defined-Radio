��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����⽸���D��6T�8�{N�/i�kf�!�6��̋"X��:�����\N(h�-����}!���1�����4�0���S��k��Xd�d���{�8�%���AHǚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>:��cG���Up�Y^����˚;���"J��+��sc��Y6�f$6�5&���z���������`dcR�+��b\�v���D���ղ:h�W��j����='�5Cq����7�r!��:l�6�Fo���_˪��k��LH�]!��0oq�1�^CO7��W�K�寿��>��h�, I���w�"�8M�@;wY�(+V��&Ns�o%�ZK�d��/��,u��y|q��g��6oD��h�5��x�+�/���Tb������Q�Q��˧�	������p��!�4�c�����oE6˞�֞��S���GWE�t>=Ѭ��y��#47p?���m�د����W,�DxjS�%	1��6ǽMX�>�M9B�Q$U��$����j�4P+����B��.d���bѢ$�wWOG�or��ӥ�^���s�N1Oʯ�衜HCk}\�>��o_ˇJy������n��)T0ؙ����*��W1�/���@E�x���H���W��;�b\*UT*Ua�.ߐ�Φ���F.���#�����T�	�H��
"a8��W��ȖΦ;1�ڨ�g'��N�"/�-�m����+�^�L��V��4G�`Y��6��Y��&x�t�[�����8e�9֎.g�A�)��"X}*_�%�VW���Ppz���g~�"�.Ru��e1�����i��ēƊO�V��k�TuB�̹�n)hx�o��+�Y��Cu��*O�����Yt�~���˕�E�sٿI�ti��N9Vp�;f@�*~�9��.�o&K��igݡ���E���f�<�f#�Æ��h41�R	k�Z(���IƮg\Ƶ�[�{9އ��sbX�J6rk���Sy���k��Y�q��g)1?~��L �8b�F'��o�l	rJK�xf��������w���R�ҩf�j�����`<BUWW -��ح�2XfW�~î�	���%VX% �V� *�Kޥ�Hk�ʊ>�y���}z�H��I���Y=�������<�c�܏M����hо1QW��A?cю%�o����`��N��@��n��>Ϗ��fּ��,2�0W<����r���g�A��x$��.�e���~-N��K��d�VG'��k���S�<3"�Y�X*(R� �3� �Ս���ɜn�ML�2�Gq<���i5������/N���O��o�B��ܾ��#��c�<�̧����E@3yX�@�<��%���@�a�����W�;�����k�O1���nx�;����`>-��$���cL�h��m��F�ŉ�0�P��Q[�3���8�i�.Hύ�/KA�]��s��aT��Δ��nj�}t/:l*�>�xw���SQ��e7%g�6k ��4h*�S\������s+��	(h4��o��6{�S�#TF[ڐ)�ݻ�}40�71��8�e�g˟\Eh��q����Q�F;'q"���$!���Rߣ�o;��{0p��ؘ!��Oy��o�fes��Ȣ�_��).��C�I�]4�I� ��C���:�@�s��y�Va�0Qh��㟅Ju�4;�LkT�w;VORNܛb���^� �ւ�ㅊ*�<�*g:�\?3��I�<N*y
	I;
�=J��fD"��F*�����7-N�{ڊ���iC�=���/NJѝ�_���7�	`�%�����(�F�#fn�Z&��A"�i���9��{�z+�blw�t�<_��]#�ǀ#F�(>)�F����(�s���Ńٵʿ-Ă=�W�	�^=��S&*uU5:_��o)"{� ���/��b�:�MsQF�p_�af��N���-AA��EU�5]�c,�Cq<`'�ݙE�MzXl"�"�d?xq7���$�'�3���ېY�(���B�na�~+�핡U�Sk>��y�c5���.�M>�Y���D�M��l���~>��00�1:4q��#���"�Os���AZ�e3�q��E��1oGq
q���5��ӁB�h*s��}
c�~���=YS<����Ugd�2�j���wA,���$贜��R�/���
�W��-RdP����
�4��} W��=d��-� PZ���r6�3~c�o?38����Y�j�r="���U��}�/�>+I_F.`��1~l}k�9�l� .�cϳxά;xH9}��;K!1��s`�(J�Y�w;
��@� �˻voL.��x4ő������UE�.Y\]]:`����*~��t1�^�+{���0��:3�����q'�IP�TH�9J�W��6������g��RI�b0���޲9B�"�5��!�v��8�D����)�T�����nG� W��s�,ښ��h\�3��sј��d��4�aO������EyKO��p!�G��x�Ҏ�Cxn(A5"���&�ُD
]Y.N���S�p�����,�q�{�y��Ҩ|�G6��5����kbf�}����?�r�5 ����y��a�H�����蝶�ׂI\ߜl
q�'�V�5��3�G5����?`��'�O�M_� �VW{����Ǒ�ܦ�B6_� �[6%�i,Z�$�����PX2�iXx&'掽�o� Gx��D$��R�ɉ�u7Ni�Lf���,\T��i9	nC)d��f�H_&�w��+j$���c)͒��7����B`^��m���R�X7�Y�f�\VtvЬ���'e}��Y�W$nY{s΃�B/�;B���%�"<��;9M�`X�+4�x���%k�a�1\<Ȏ$�ث��祪	�]�/��I�=���F7)���FK㢬NJ<�t�.��'_�Ċ��{���ޞq�y�M陷�^��#��4�ђe�'�s� 9�S�f(H�l7�1��LC�}g�e�da�lÄ�K<[��r]2z{M�l����u%�(W�6ܛ��5.Ua��.���,B����*
R�â'}�'ðz�7�I�e�ř_����[�OPT�l�r�y�(�U��9�4}-���S�>�>#������&����:=��Iq��vT���Y����r��Ť�I��lH�Pu
ލWܧ�;�J�u�`��~���G�SI�o(��W%��/�P�K�0V�q>�L��K|�I2��HA�#�ѝڀ����=ASF�K���_��<8�)=�r,�u�J1Ç��S	=�5-��0"����1�{>xe�$+��sZ]{[qC1�*{e���O��~�<�b>f�L7۶qG�� N��I�C����A]>�Jmh�w!z����1���>��5-���LV=��3���e���^�*�C���#����v�2m��;u���O^��5/ Xܩ$�l+�"���/ZF��O҆Q�9d�����ܻ#��-���)$��~
 V	st��5�u��؁��S��;�e�|N��X,ye3z<��摂��t�Z:���K�9��CC�V�<��щ �2��tE<����c8��6L���jВT���o��7No&؍�>�b� �A��zI���MF�޽"��Ru�5/H�_�W��]k�t9���</�>�4������d07|i5���K2��Wr��f�r���L�d�`& (R+�n4R�r�����RIJKF�ʨ����j��Q`�F����o�~��k� �u��!f�Z}+e\f�
J 4�c$&qa3&�_ym�Xs@���y�$WW�G4�2�疐��Y��M`���Qm/E\�2�K���������?�ul^G�w0�e��T�=�O� a�8���[j��C�g[B��FpTZ&��k�w���{���c�����*(е����p���ժz��V C6�=X|,�vr���l
����wl��m	ENX��ѭ�3���т+_��K�3N�� K0��"2LE�7i( v�s<�����鱁Rȇ����5P��⿶vN��E����[�n
,j��8!�'3+ ��Y����	�8��oQ�A?D��~Yَ����ڿ3����jՄb:�^2҂d�+ ��4Vְk^��^�>A\c�Y#����R��S��N{NǞ�m�4���Zr���ӝY9Ҟ&���& ��v�Q{�dW���N�� '��S%�F!L�&��]�2���Z3�<leeϡ�)� �
I���S�5��D�b�IM�L��0M!�蟨W��2�gI��,J��2"@"���4g�-��
/�bb[��c*h�o�'��x�"�ntz,�|��kʞ 
�EG_�ʓeJ�8bUO��"MWLp�k�"mvSJ9\b�����멳[� �H��ͨ�����G���T�{�e��4���t��T���sa%d1�Ed*+?椺/�2�mؑ4��}ށS�4���L-�^Q����Z�#�D���������OZd�-䫫��m�IH��*�,~)��+��v�W�3�:�~�]02��Y�	�K�d?����Ҕe���U
�-���l��E�e���J�W�%ӵ���d��k���K�@�lp��8�?� j��Ǫ"�mW
h�/����*�L���
ٙ+�kE
傴����� �[0f�ϖeB����ۑ����ـ�ǧ���wU�:>��q�m��&x�D����+a�����NC����jTd�3X�|
�n���X��u�7���P���cl*�ȧ����mLk��$��?sH�g��P$�o@�ħ=�t�,�f})������d���� �#HQ% ��[�=�){�T�}���r��@��E�>Ńٗ\�v��x �M��п͐@�W TI�}B����z��*��dr�Q�U�������aV�YC�F�+?���o�����Q>sm��뮦!��_�cb�y3��
��2���L�~�Y3b,�B�\wZ7��`�u���G>D�yd���0T���Uu(-�y�3(�w��Y�p၆̯����Ft.g>��^�4�Ź�[��U���	��lDM��3B
%�=G��%-4Z�|���q>g�Ȼo�r0�lj������v�&����M6��|n�����zЂ
��A\	q��0ד��ۍ|S� �x!Ѕ�~�SC.*h�����p|�_UeÆ�4�[�"1p�K�ĩ�j.=� éN�,u)2g�M%70�r\]I�N2�t#�`DS"�/�����hY�Z�)���`�pt�8�FM�P[�.�M�a��H����Ob���IˑaӞh�`�dp�J	�ܺH�ेg��)�� Q���:�n`h�M��n����uZ[��y1d@�qYL�h>�몏���V��o�a�
SLe3��y�HJ*�+�4i9�'�Z�������8�wH��H2����E4eȇ{�%;Ŏ���pS_�.��6�����T����&>��eJ�䂠t�ĽS3�T�S��`o#��Pл��Kv�+��c��d�x�7��:-IB���>�=i�>�ֿo��5�N�5C��im��Ӏ��\��NC���z�vL�*B�еET��(2�b�u!rBfɻQ��Q�_�
XU=�lz4@� �4\�^ةh���r��2���$#���
��0����=�p���2Z��u�_��7#R�8���;]�A��UR�(��Z
GXve��� d�0��7w��Y_;�����J��&ʾ*�5ݍ�W���V��׬2�	o�1������z~o}-�p�*GZF�,�#j{��M>�r�;�d�����ԛ��YO��Q�¿��{��#v�&�_"��4���"W^����F���ê��H�\P�<���7J��m�wiMJ|��pK}���
�v��n����|�3���
v�H:�Lͧ��S�����Q�k�~X��	q����b���f���������?��9�`���s*��\8�yI��q�i� "��zz�GɐB�B��:���g�~5s7]Hb�>�'ऊ�/�SN�ۇ�~f*����ۖPӚx�(��_E;�(�0�Av�Q7�7ȪMjt
3�H]��!�贮��L�C=�K�F5C�8Hj�2�?c��F�ۜ�Ǌ�R���73�IE�d���;�/ʟ�����t�����!�I#Fy;b�a����o �CF�ǁ�Wv�2��]"?w� ��a.JPa�.]ep|�ɠ2d���j)�%�sp3:[v�T����K�|��.6jR>��p���z�k���\d}{� ����4�8*X�����zL7)��i6�ud����Ln�˅A�ڊ�14�Ώ�r�$c�gT���8xۥP%ąr���].�K�l�Y�9�C��E6�#)|�v<�ڤV��@ �jIh���cj�;>o�)����$�WfzU[{M�1>�2e�\��R������g���8�d�k4,*TJn�57�4�s6KbݶP4�^���J3��g%m���