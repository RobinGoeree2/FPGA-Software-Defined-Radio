��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���G�H�ƻ	�"�iQ�����3�7Q��㼫F|�ݽ0��@h ���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�s8�R�	�}����T�l䮱}��V�W��]��;�Iώx�t���E�L#uc��WŬ�+�-ޗ(huUPh2�ⴓ������g�ך��_�L���$�1�2m��+�<4��ˌ�ň��h������R��t�  ",�N<��;��� B]�pE���	x]̃Dj#^Da����M���Af\O��x^Q\7�z����)�,�˛D��w���旴4�����<��a��rl�ʩ{�Bf��Sd,�ϱ����@N1�w�0XL��t:w�~�gm��+��9��kT!����Y�f��a�Z��VRX�U�~^MZ��6$%*Ѣ�?�.��l	���./����C��c�S+d?S�7�$�>��8��{9�dcCY�=\O�phpA�J����L�=l�)��%�0|]<w:�dh��0�l_Ǒ��\洽<�p����=WL����_U0ϣ�2$6�sIMǓߥ)��ཡ��!�`�(i3!�`�(i3�d �^�z'��� a�~�d��W񳳢�l�"��!�`�(i3��M��)��ہ��-��8<�|�(�#��_�1��k��5@��7���[l�A̱F�9�����Fz�!�`�(i3!�`�(i3��T��� ��$�Tnf4w���f\P�z��8�8���"zɰ+�*IZ5AzO�  ���Fz�!�`�(i3!�`�(i3*���C^��#W��xW�tI����h�;Y�R��㕞o7 ��r�g���DD6I�a�W�t�lE�f���p!!v*!�����ӹbm�@���*�n2�=�zOc�.[K��m�:8��(HE�����!�`�(i3!�`�(i3>[�ݗ*ͬC�g.jq,�W��E$��"����!c�����=6Ws��$�Z�����c�sȸ�"rR!�`�(i3�?�W/)Gdq��c�冭B2,�Wpv͔���Ef���=R�?��nQ�-�j��Ő!�`�(i3!�`�(i3������!���C�/�y2+Uv�_?�#׷�`�:\�t�Z�f��r]+q��p4/j��ㅑl��o�ڭ�������lI�@�$��$��5ف�*���J�]�]��X�p0��o�_Y)'\y��=�2�!�`�(i3!�`�(i3�K�Ǔ�\�h:qP�
]���J��:�I,�D�y:#9�]�B�-����;���=���0)�Myիnň��h����]ߺ�`@�Ny.��d�7pp��8X�˞�DG!�`�(i3!�`�(i3p{���gM�k���lh�&ĵ�	ƹqE_���RQ�
�)T^�b�k�@����S��l��ׇӭ��!�`�(i3!�`�(i3��sƲ����e:��x����7>�����D/͘B���&,��*`O�4��.�V6���{ֱ@�,z���h���iI����p264!�`�(i3!�`�(i30tYK�yPVq�|`kK��I�+�:钾Ci5���y2�����J՝�K�y؄@�!�`�(i3!�`�(i3+���6>�2'5�sZw��Q�둩��n,��'�\�n�~��q"P�H�oe��C��c�S+d�J�Г��f�u�����!$檦!�*��Q�`��=vݖ6�F!�`�(i3!�`�(i3�s�cn0�u�A�qL��D24N<I8����\.W~C*B Ɣ��(J�f�w/�BWSl�p}�!?��~�7����*H:Ky}�	� �H��*%��6�A:&�����R�<���"n���X���K�y؄@�!�`�(i3!�`�(i3����ZY��@������'aM�Q'��R���?�:�_"����kYZj*��$	�5��Y;ab95c��!�`�(i3!�`�(i3
�;i%?j�#ʘ�s�V��R��x����'�;W���U�WN�b�D�#��Q4�����Fz�!�`�(i3!�`�(i3�j_xK4M�gҞ��Z_��=WO�V2y/�xe��[!���+��iDM�����sȸ�"rR!�`�(i3�����$��뵮�a��K,<o���,ĺQ=X�5�I��Pm��G��ZZ��PY�ׯ
`�!�`�(i3!�`�(i3%"b��4P#
QjK��18*��#�N68��_kCڔ��&���D��L���_�L�����J]5+a�#�$�@%���Q� ���6��H4�
� �AH��,�2�K��0ӵ鏽�闇�{_������ѕ����AcX�pA�o%����RL�a)3���ʉ�N	:.���n�O��w��)�R�1z!,!�zg�Z�$��,2�v����"�D��S��<������k�bv��;6�ThI^����7&��N��K�r?���\z-��EM���
+����rx�]�V��\#O���o�x��`�|>���P��f�>�٘\ׇӭ�ѯ��[���g����=�E����F���8�TP֪zw�&��Rb��Y�W��OC��E�}��W�p$ܢ��{&��ؽ7$�	�s}��[�X^#��˄��4X%�_p<s/'^@���`���a�ٜ췽��/���ʛQ�REzv��wvC���		�:���ʖi5	�ݐ���E��?ؚ�v�}�h��g�I5���S��$�m;8C��<(���}0xH�����PZ����M=�_�mD�ʮ��SJ,8��µ���x�_����eM��Ų^Ε���}�P�������pC-��h��☂/x+��s(a�L�"�,�9�{��2$6�sI�حЄSZ�h�5L��p
� �AH���g���	� �b5z���lR����W.=�2����QE���Ý�M���AQ �����Jw�)��e�0
A���l6��n�'F�H�(�/�r8@��Ƥ2���_�xm7��(С�"pX�����U�?��+�x�8�n����Oq:m�j�{_5Jwʛ���[E�8z���U ��?��k�Jd����r�>>7�*���/���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�tw:g�V|�hi��p�7��Z鎬�����R�LM��ħƿ�9c�5(��}���SaB:��}������<׏^��|S۸�Qk�� h����|H�<�'��I��"ˍ,�ʓ��M�%��Qe��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcd��q�G�+��T���jB�Fg�Y씤`��px��.��r�M$�*� ��]���t�iZ]XF�������̚ԅ1Qr������i��E����F���8�TP� �B�ݿmŞ�����ȧ���(�w�D��y.�2ӿx<�!�`�(i3-r��|ڑv1���ȵPʶ=������Y�n=n�k-�;��H`��!зq8�ЈR���b�>���4�ʛ9�0�̳���i�#fC/�����Ul@�;��Q.�KUfc�^~W�BJ9�c��N�w�t�Z�f��=��9�JHn��z����A3�lz���+�8ΒՎ h.\���Z�
�B�qA����ܱ�y�s���z���+�8$�ݛ5�CN��������+�J������܌��14�:v~E�)d,�vd���x����n,��>]��e�
����n�4];ˍH����_�.C (��o�e5�3ͯ����OtB-r��|ڑv1���ȵPʶ=���k<��`���@���[K����Z�ą��v1���ȵPʶ=������b��˝Sz��E�4.@��n̈́�����9�3�{z�k�/���i� � �	{��Y��
�iCY%T��BPS�)37J*u>����C��U���e�N�By3��<Z鎬����A��:6])����7�RWk�bU��e��I:gϔ�&��s���q7Ê7�E�4'���Xw�,bxqX�a���C154�EY�o\�J������m�F�䢝{l�f|�ό���.ӽ����
�Pm����ҋX����>��l%i�-'�b-����׿�߼�E�]�!����M[��ǢF�\�h�7Ê7�E�4'���Xw�,bxqX�)����p��P��OfyN�D�li�.���cQ>N��g������cQ>��� qv��s'��;ɩ��}�t�*-u;G�w�8�}?��]�!��	Ǹ�y85�C��H�����t�Z�f����8���D24N<I8����\.WS�UE^��\�HP@�a%=dϖ�i�q㧵�0������0��D��L���_�L�����J]5+a�#�$�@%G���V$��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h}|��XH��9��p#�7ڜ¸<�X��/~.)��3\�R�F*}�c}��uOA�ٗ��J�"�却G�G���cU�J;��	�yE�Ss�x-��A%X�z²���ʓ�*Aj�I�e���_�$��*�yW��Xi9�
�іm��U'�k���W�f����ހ�Fhʢ!�5��=l�U�-��#x�۾����!d�h��<�qƂ�$�������i��O��$��Xo��ߌ;޴@�,ԯ���gn"G�q�������b�3!^�3�@ym�-f:2�	�^����Ћ�l�Tq��W-q�C<{�uig����V�dN�<@Iv�O�ȕi�l=I��nȑl�5��̄qbqlФ�vt�q��gbb˸xZ鎬�������(����\\�*�}!�X�V0Up�rP��O%�ud]�M��+x�r����l�©�]t��):�Z鎬�������(����N=�[��e���ZF��ֱ�q������m�q��|�1��TZ@�6��7�){`4�2N��n�`�*�������r���Y�{'%s�6F���y�b.�hFd=��¾ȼ�u{*�C<�3�@ym���Ζ��1tSjv��37y���� ���30��w�w:�;�jmT�#,��T�����\_���/]�l�����&G�q�9�ͭe���PO�my$�N�����'�ډRa])n#���r������vf�<�R�{_8�Y���0�-��Q����ƾ�x�\oqv !�`�(i3yY2�̾���U�;��tS�$bnNfĉ>99��A0ok��[p�#�_ wgf*��$�Q�����S8�&u�η��.�[�X��=�gw�⽒���n�����:=�e�)�ή@���P��� �Uj�.�B��0�9�@�`���}Dq�f�Goj ��6^�h����!�`�(i3pı��0����%�m1%�Z��3��w��\�W�ƍ2���lĵݓ�W����l3]�T4�0 L?ஹ�%�ԟ����U��ݚ�Н�(*�O�q�ͯ�*�d�[}�N�`2���K����A0��s!�`�(i3�u�24��&~e�e��E{��h5���՜����|e"ʁ���MյX쯢86�	Ղ�I8�y\��S��z���wb��Z2!�`�(i3U /숇�]�	bC��<-�;S5b	��T�.�w؀�CF��6��� m�#;[��U젩`#FW8�	����C��s;��}Dq�f�G�&ց�*�=��
��P�n���}���S.�3��"Uʡne�!�`�(i3pı��0��Y�]�q��c�Z��3��w��\�W��@�����ݓ�W���D��!~�4�0 L?ஹ�%���EXc=Sq�ݚ�Н�(*�O�qm͈���߀[}�N�`2���K��m���
`��!�`�(i34r2p�jg�&~e�e��E{��h��^9�Ƣ���|e"ʁ���Mյ)n�B�D�	Ղ�I8�y\��S��z������'�!�`�(i3U /숇������<-�;S5b	��T�.m�P��/A��6���r��(d��U젩`#FW8�	��2g���ܐ��}Dq�f�G�&ց�*�la�T�H�n���}���S.�3��7�E!�[!�`�(i3 |������if��Y��Z��3��w��\�W�ed�N�-�ݓ�W���	�N�M���q�嘝��ஹ�%��2V[���X��ݚ�Н�AL(�z������0`�?�JY�)�q��ڍ�����a�"��6���@�HN��R���ء�I��$�S�in�Ye�ήT�C�5y��;�@����gGɑ1tc5+�o���B���+�J��P/;D����L�E�$����Y�Q w�)/�L�He�-�c,!3�?4���R;7s�9���o�jƓ�[����ըi:�HCaIMl��*�>^&9@^7&ģM�I,�D�y:#9�]�B���' ��Cҷ��ecx�S�����S8���IO,���������9b�S� 7�v�ԯ��Q[R�7����n9�O�M:R	�d2}�#�l�1����?����pҋ{y����x��F�U| c�]h��\
�QQK:2i�ȕ���Q��i7N�_�wDo�h�'�t�Z�f�}��+��\��5��,bXh��d���!iEOJ�uxm�PQ%cp��g%`5D(��A0�r�P{��Lג�Q^�MY:�6���;b��g��U-�e��:���j�D24N<I8����\.W��/z*x�n;��|B`q�a�i��E2�DZ�⸖�A�{ �I��/|��6M�Y4E&�|=��s��$�Z;��|B�8��w@<;0V5����[�b���^PQf��і!�UDl�V��b)N�u����S���╔�V�T�99�M�g������E/��F��An�D�	+���G����?����2�T�$㥓�@qO��Q�rG�LN_�#<���ӟ@^9�C�{a�?Ӯ��A0�rR밉_@UB���_�w�~��}e����"����׶h���G��w�L�IX0F�MV�ҁGGSoJ̈��:scX{�X!,!�Y��B
��v{�*�g!�`�(i3$H#Ö涅3�<_�ټ�G��z6!��TޅiL݃g{~�5H:csK�g��$�Z��cp6Dq��;���EWrqi}�Еi!�`�(i3���#] �����a���'���_�)��Ƒ�^�2�"�,�>E��ʆ�In��t�1β��cp6Dq��;���EWr
Cj�R[z�����/�jݭ�F����=@'ѥ��~�26��\�́�T[)�W�=�k�l0��F��j-"{b����$�Qu�84�^\���C9*�¢ڲ��+�J��&�3�Ck%̷��q� �#�� �\�7>�����ǚr��y�h'( Ik\D�P�E6����{���$�Qu�N�#f���C9*�¢ړN5Χ��F�,ؚ��XJbk-����'�\�n��6��	���`y���cp6Dq��;���EWr��Ϗ�2�l~ޖ���[�ć���7)��]&��:0!�~�26��\��C���u�ÅǷ>���'hZ*rw�w����Jjz�O.C��|#HK���d��JXl'�T��~��Uг�|<!�`�(i3���7�
�Q����>���>:Y�<�!�`�(i31}�ั):9��tf��!�C�U���T9� )� �a;��d8Q�X놱�/Q����!F�G����b���/r�P!�c	{�}�|�sT����%"��/8�NJhd��
���G��RVf�I>A\!w��Ip�9�O��F�`,9�H�W�I,�D�y:#9�]�B�_��wBW�MM
��,=*A&-�Ri!�`�(i3E��\�����۪%Nb��B�i��@�7FB �^���b��n1��$�1#Q��e�.�:5A��pfĉ>99��R�V�"�0�!�`�(i3�j����D_���w�]Jq��BѲ�+���L>!�`�(i3%0Z�M��L��՜-)����&}0�@��}Dq�f���Ě�����}Dq�f�$L��ǚ�ė�v|����Ƒ�^�2��T�TN��<�6�Q=�k��M�1}�ั):9��tf��!����WBe���	IB�_k�e�8��B�:5A��p���F1������$����sR�I�uS+����:5A��p� ͷ�	��@.�$�_�`
 ֢��؜J��v�W�Hl����A�T��K�P��-j,�`
 ֢��؜J��v�"֡�7�=�o�l������[<�6�Q=k�oR2����f������F1������$�����̪S�?P�|���������"���Ȋ�?ӳ4�;Ⓠޕ;j�j�������"�
�T�r�5���@dr�����S>�;�u��tF�{F#����]���o�ݚ�Н�6S� �*�����$����sR�I�uS+����:5A��po2p��8§�F�^�S�!�`�(i3�JO�'��+��K�L◁���*�8Ğ�
ҳ�͜�}Dq�f�1}�ั):9��tf��!��Ϗ�2�ed4���Ȝ�}Dq�f��1Ƈ��,��v�������Ȋ�?ӳ4�;Ⓠ�X/�7�D(��{���>��%��u����Ȋ�?ӳ4�;Ⓠޕ;j�j�������"�
�T�r�5��� л����}�pd=!�`�(i3�JO�'��+��K�L◁���*�8A���B
ԧ!�`�(i3�JO�'��`gw�T�с֜>�E�2w�f�%!�`�(i3Cݮ2����yg�^�a�ݚ�Н��i7N�_�wDo�h�'�t�Z�f�t���p,�7�g��U-�egt�n���!�`�(i3�,}უY�1��� �U��֜��3Vr�O���J�\���=-�aT����-�]�l��O���0�J;���[�uV?��?s�ʭB�?�`u��r��!�`�(i3z���r#� ?����6	�T��u~��t����>PQ%cp��g�H���~��!�`�(i3E��\�����45��"���G��#!�`�(i3��i��:q��7>�����ǚr��y�%�!��U]�ߍ�2d��3џ1�F�Z	��c*�n9i��g��It\$�ݛ5�CNc*�n9ie�{�W!�`�(i3�8@�MUn�=x�mdE�����o��26h�W�5��|���}Dq�f�`
 ֢��؜J��v�S1��6�uE9�+��՝� s�#�K4ZRP�����9�p:}�L���)	�8VڂK�ykv!�`�(i3@?d�s�8K)�W�=�k�Ҟ�#�>��(�%���]v1�_ُE2�DZ��[Z��.�~!�`�(i3a3@��[/�L��O��pXJԱы!Te�g�`�f�ݚ�Н��̢k����J�\���=��}���*rcxm�N�e�{�W!�`�(i3�uz�#-]iyQ���4��}�@���_rS�b�8Z�AԢ�a\蟘�26h�W�5��|��:5A��p��6������S>�P���b�g�W����C�M��!�`�(i3�5ߧE4��!�`�(i31}�ั):9��tf��!��Ϗ�2�ed4���Ȝ�}Dq�f��u��A�0���򴶽!a3@��[/�-=�f��W|N�Y������f��`ȱ���}Dq�f��5ߧE4��HN��R���IX0F�M��)��ֻ�aD�sD�.�g3Zv���� j��LY޺���5�IcV�s�u��6h�����T�ǚ�=2�L-���;@�1���C9*�¢ڵx�xx=�K�+b�&烈�|����b���0��Ah����+x�r�}�9�P:��&sq�?��I"�,�>E���2,��T���$�Qu�)�˥D@���D0�y黛}�)��/oq��WX ��b�FP&s��K���!�`�(i3�a�\�����fZ���o ��b�FP&g�P7�#�!�`�(i3�a�\�����fZ���o ��b�FP&;Ε^���N>I��WJ��a�\�����fZ���o ��b�FP&P"G�wk�\����b9���1]�?��� ��b�FP&��㟷7��!�`�(i37�ܥ��2�'k��� �&�C�|检+�9�jɲ�1��� ����P�7� 1�ж� �4���܂��+x�r�u�#��nt5޵3{�aP"�,�>E���Ԗ/�����IO,��������;�¬pX��g��U-�e�,���6+� ��b�FP&|��^���#	#vqG!u<�a�\����N'�D���h��㉊���;���EWrr���ӓ7l~ޖ���[�ć��@�|��D/�O��1�(&�L����^a�nu4Bޗ��jw�	���;b�-�2��⅚ld��b�M�⅚ld�^�R��m�|#HK������ �'����u��r���@�d�u�G_"�|�2�d��-��!�I`��G��T'����ð��T�ݚ�Н���=�g�żפ	�?9Pjp������PN��7�v�ԯA��bu�x��ݚ�Н��H����˜�?�������gHucP��#��s�gU-W!�`�(i3���	.Z뵫S�"B؟�r����ڵ���[�m4Z�N���{��c�C3M�6��A*�6
�7!�`�(i3�([��B�{?a� ~>>ը܅%Gb���U��w�1tSjv�!�`�(i3���F1������$��ʆ�In��t��(��+�⅚ld{ϝ�[�{!�`�(i3���Ȋ�?ӳ4�;Ⓠ��c#�Խ�������"�
�T�r�5�!�`�(i3���F��O��ݚ�Н��H����Jbk-����'�\�n1���R��뷅Kn�;F�Q��s,�~TM�e�w�Gr͍��Y�1E�c��>ݎ�T���r͍��Y�1� �54�T!�`�(i3�$�#{dC�(��mp���Z�{/J���#D}(��26h�W�5��|��:5A��p!�`�(i3E��\�����45��"���G��#!�`�(i3�̢k���!r}<ﷹ�Q^�MY:T1�Ɓj9��jg����ΒՎ h.\���Z�
,�/>��a���9w��d���[�,�/>��a�r���m�5��ݚ�Н��0�9&،��)���4�����wb���H�1����?��&l�p�q,!!�`�(i3a3@��[/�L��O��pt��1#��
��}Dq�f�՝� s�#�K4ZRP�����9�p:}�L���)	�8VڂK�ykv!�`�(i3����&��vL n9-�N*��D�x���Q���kO��u�:�HCaIMl�i;��B��}Dq�f�!�`�(i3�JO�'��Z�UT'�vL n9-�N
�T�r�5�!�`�(i3\OW�:�ݎ�T��߶Seͪ��Y{Y����H�����1tSjv�!�`�(i3�uz�#-]iyQ���4��}�@���_rS�b�8Z�AԢ�a\蟘�26h�W�5��|��:5A��p!�`�(i3E��\�����7}#�ouߗN���g�3$�J�5'!�`�(i3HN��R��bP�63Z�t!�`�(i3%ʴ�ɒ�L��C�/�y|2I��js��'Q�:�H�RtV�^!�`�(i3{[�ב�C���#�'4v~9��c�	?�N����!�`�(i3�����!�`�(i3�H����y�A�룘8�u?��I���y��lD�\K#|�t�}���zd�Gͦ�Ũ�i�/v�ы�����!�`�(i3a3@��[/�L��O��p8�#.��#�C����!�����!�`�(i3fĉ>99��A0ok��!�`�(i3���F��O��ݚ�Н����W0�]��e|)0����n�=�H����ʒ���)0�x����VY�+��I�j� �&u��r��!�`�(i3{[�ב�C���#�'4v~9��c�	?�N����!�`�(i3�5ߧE4��!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN��Ě���aT��3G�IX0F�MA�ٗ��J��i r�_���(=)7q�'GWy�I]�o��_�Rv�䩲$����#��i��ȭ��J�E�b#�T_0����k���,� ��b�FP&s��K���i3<�f�D.`�Z���N}�m��{�K|��S��Z�:i.ߋg���~�26��\�v�F#�5�f
���K�����o0H1��M.��jJ3�9�C�s�4d�G}%����3f�Ɲ�c�M�%K����`�7�癆cgR������������ h�ҩ�Juv��D1�|�F��>�X6�j~H�RtV�^J�N�d�	4��'�����R�Б΀��E�b#���P��0	J2L0�jdc�#����nS���4W��C��#�a�ĄqcCl���<jJ3�P�}#���u��r��y��j��k	y��C!��AVt���!ɉO hdU�lP�k*$LA(k��'?"�5�_Ym$�T9w�[:��q�HN��R��bP�63Z�t��Ě���!��"� +}0�ʂ�j�Ï��	�l�lM�3 H�RtV�^d)ɓ\©K�Śޫ�#Wx�Ա�%��ݚ�Н�:
��x�{�\��N�Ś�-����!�`�(i3����i��dq���f�e���v[v%��?����9<���H1tSjv�!�`�(i3�-(�̿x����VY�+��I�8��5��_� h�ҩ�!�`�(i3���W��Ȑi�X!�!D��(J�f�"��3���!�{K5~�{ӭ��J4h�!�`�(i3f���Ն� ��%�D�v�l�Ū�TD���7��y%%9���.:��Q?M8�f2!�`�(i3�wbk�$q6��@�h��q�hgvCq_c�!
�T�r�5�!�`�(i3>�������G��#fT�R�7h������e�d��I$EI[��(��!�`�(i3!�`�(i3a�/�	5�5�V{��RCJ�����@�ĵm�ݚ�Н�!�`�(i3�?�JY�)�q��ڍ!�`�(i3����a�~9��tf��!.G�9^&���}Dq�f�!�`�(i3�0\� ��+s��K���z�3�0�M�E���U�6�'�)�Բc1����?���U�	e �!�`�(i3!�`�(i3f퀔�����̹�d.ň��h��:����E�c��ދ�+%C�@�&B��l��row�	�r1���4i�'�n��� �Ξ[�s��\2��T���W?r�Q�^8�bL�1p/-��N�]|-���"�s������f�ʯ�`�D�ʆ�In��tN��H3�dv�c-��?���$73�!	�Ø�e�!�`�(i3���%>�rG40�RS���$
�)!�`�(i3�����!�`�(i3�� л���I�+�'�=�o�l�9��V�9!�`�(i3a�/�	5�5�V{��RCJ�����@�ĵm�ݚ�Н���6��w=\��*ȜD���|�]�)�Z����J�]�]K����J��!�`�(i3!�`�(i3a�/�	5�5�V{��RCJ�����@�ĵm�ݚ�Н�
�:qEpCt�w#��@�ݚ�Н�9�O��F�`,9�H�W�I,�D�y:#9�]�B�_��wBW�MM
��,=*A&-�Ri!�`�(i3.��J�޺��:p~	E�<l��uE9�+��!�`�(i3�d��R�;Fc/�p@�dB<4RW��rS�b�8Z��W�6?��O�M:R	������f퀔�����̹�d.ň��h��:����E�c��ދ�+%C�@�&B��l��row�	�r1���4i�'�n��� �Ξ[�s��\2��T���W?r�Q�^8�bL�1p/-��N�]|-���"�s������f�ʯ�`�D�ʆ�In��tN��H3�dv�c-��?���$73�!	�Ø�e�!�`�(i3���%>�rG40�RS���$
�)!�`�(i3��Ě�����}Dq�f�HN��R��bP�63Z�tHN��R��bP�63Z�t��Ě����E�i�m}6O�D mWN��ܐ�}ĢƝ�c�M�%K����`�I~m��DL~΄gO�3��|��[���Αo��p2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc*?��J((