��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����⽸���D��6T�8�{N�/i�kf�!�6��̋"X��:�����\N(h�-����}!���1�����4�0���S��k��Xd�d���{�8�%���AHǚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>c��mW���rJ(���/	���~J`2F�x���4W�0V�y��l]��X���8D�G$�ۻ��c��rk�E8o��W��z�����O�Q�F��?-_�䰹��Ny����o��:���l�,�:^�G���G��ta�`����k�?W�lo��]/ޫ���PȚ�-�sx��l'��
�lX�ۦ����.�v�D=�~�4C��~�h��6$�^�;d��G�M���Ѵ�S���ګ�\�̿��*p?���/(�D�"m�Ƕ?�I��ɑ�[��r~���}��5�Y-ݮ�j0��6��<��{=�����A_�}Q3�����mA�ܹ�!�Z�^G�(�v�P�}w�u�4��Z�!W��o9F� ��]�xh��h��X�����b���B������^'��?��[S��]������F�אo\�:�|�=���h�L9MOB'"�:�8��;c�702��cҐ4�%��N8�~	�C֐���ef"{��F#��6I؄�Rmj0��)x'&�)@�A��� |fӤ@������H�<��]��G	]N�S_v&=[\߈wH�T�HG1 Tv�#�E�X���?���ߚ�6�O��ĺl�9ŋh��d�r$P�Xb��*�!�s""��6��z�����l>Z�U�~�]'@�M�������	Oc��#Ue���(�wP���o�E��,�C�5�� :����j;^�����ِm��[R��;{P�x�2����m�ix�Ͻk�}��4��q:N��?�3�JU5����ۥ�J*���ǈ��w��Z}A,����Ӂ���8��6�2!
�E7ѫI�����(/��$1�`�x,ܛ�zO�eM�G�hy;|9u����*����k��3����/���SC�/7C�r8�����兠�#3ȥ^���=�L94�Y�V��P��7�e�Ç�-��<��3��a$��"���O���b}	CSH�bbԱ����P�j���2��Z�N�*��'��A����!�������($U63>��� ��U�r��BSN�s�5� �qͣ'�w�f*���r�H���<��W�iߖ��N�Z���~j��z�RsF�x��XI�0e)�6d��x��򹀖�\�	+o>Ҥ>Q��p��(�e�բP4hɰ�@
��U��XNeq]�?�K����k��ͷ6���G�>H(m{�H��KC�����!����鐸�o�[�-CU��G���!h��e���8�+�>(&c(�.�o,on����Ya��@.�d	1'�jƻG�G�����/�����E���k��m� �O�1������X��zDpk+�&�v]�NN�%�D�5R&�F1�Զ�Za� �l~��>ss:��el���IR��d���g��֋T��ϔ�i�}����G����i-p!����t�q�.�S)�W�;v���D�Zӻ�h��v5����3P��!����'�]��
Rm�|�?�%�R{�W��-�������++���9)���$&/��b\��$\�j�Q�u*�~¡���}m��\�=Z0��с� �*�x�M�>ّ�Dy�y�5m�V���
&�R�`�In�\�Z��ÙU��^�=�U���fM�Ŕ,e+�\^ĝ\������'5Ah^�+O(D�1 �u���PW ���q��)~�{%��?x<�,�f|)G=���2P1�;��y��A.]����:hF�(X��<��ŴV2��b҆��Վj}��<��(�0�TϙS:)d��o�*�4e�*������f�g\�|}��Z����{�U�v�7��)?[�pnr���C��`UJӾs��Y�� K�"F�/��h����}�Ij�%���[h�i2��z��W����z蛵��b&�:����A93��7�j�|��~޴�x�Ey?�לT�:����f�������N��p����F[x䚔�G��S��K��f�X���b�v)��R���tL�����ћ0� ��(����ZW�.	���"� o�ĵ-xu'[��2��/*,dfl���h���MT���~燌չ���>�kdK-�x"��L%s���5��*��gn"��'��t�)�OC��:W��vU��D�~J��M��<"�b���G�ۏ��ѣc?�0PB&=h<�y�������/hxī���4����B{�	�B��}�A�)!̼弘b�;p��i_�@����F3<�]�X��Ǯ^(�Ά��k�7�URhRԔY�2hD@��֛8��*�3M��?�S8\(� :�VW�� u���uI�}�o+n�@SQ�ܙ�/W���`a��m�c������A6z��fG�!�?��Z��Z�W���g�V�������(&!NV�� -u,��rB�R�+��n��) R&���Dn}���T�����Jö,y̓،~������<�+�Z�����{�����&���A��|��;*�g�U0�Z������r�JL"M ����-4��p���!�L�ґX���}�m�����G�G�*���SJQ�(jb����< J�0��ڶ���C'�jn����}&l��*�U@4�w��-�1?�X�m����7���]�b�%=.���ͻD���^��'�1]����ĹP���U�:�axlB���S*�YC��{��o[ �.�_V��Y!���0�+���?H�RG�Y�w���g��0���(�m`LYiR�];6���~�����
xBfR��'Lk�[��"I�QBC�&_�>ˋ��3ӓ��s�F�_r�,y������&ۼ��|����`�j����'��r�D�ӵ��U��@ng3y��8̨��4j�ߢ�j.��ʬm���N"�ӱvH�32(W͉��FJ�;��c�,�����ZI��Wk�6��_��S�}ߡͱ4�m�����`uJ0�Fj�>�F�$�ډ
�!N���Ja�WR"AI.��d��aҹ��JI��	�O��{�4'�M\�YI�I�䃑�S�g��b��s��ǥJ�d1z��^d$�b]#�V.GR1!��kk@AJҨz�ULr�h�?����sn�ۋm���g6�a�(���o���*�"�Zۼ��õG`D_�4��x�o��!8
�O�U�������i^˳A��-�.�+.d>P��g H���N=4�\_�C�iϠŏ�iH-Jh��|ͪ$p:#��k�p�N�m5��6Q�u �����Y�}|h޾"���%�FF��H���0�]Ϭ�d��ĉ�DA���AX
ϓ��6����^��x�礿ͽ�l���(�����0����M�Ƃ��g�^Q L�U���
v`l��$