��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����⽸���D��6T�8�{N�/i�kf�!�6��̋"X��:�����\N(h�-����}!���1�����4�0���S��k��Xd�d���{�8�%���AHǚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv ��i��X��s�-�Q?F�`Y�������� I֏�׋������H[��9����ۍ: ؕ��6ж���Q��" ��y&���Y	6_���.���M�ݟ����k����
۷j	���`a�s�Yot1H���\��b��x(5�;Ƈ��ܪi�d����/��%:�q��P���!Od^�_�aD|���RE��3.y�v\5UZ�d^�?�1�p�H�c��ZE���ǎ,�9�`Eb��K��B'����\f��Y��p�}�t�ra� �_�wy)i~��*;Yh�tn]�:�H�z�{E����Ji��4o�CL����S����ȱä)lSݫ��op�u�����w2dU���OMv]�L6��Rn@j�>p�r@P`������F�ZI�������6��;�}\ʾm������xN%��_����m($��JO���+H�B�7;��pְ�V�9'������R(���8����(p�/.��s$ �Ȗ��A����J �A��[K�p�lU��+2��������oˣ��mzK����>�~[Y���܆��2y� �5��5Y5Z5Up�����sdҙ�IX�	߾V��|{��Z��
h����}S}Q��H��K"��nb�`�.�Z���f�fj��c=J|�I����&�w�X�r�\�®�˯�`�sP��B�������f�_��	��8��\L,�1f�.};���e)w�����d�ٓ��ksn���΢5�IL�O2��m,�����2O��WD�%fL���}Y�"�jb�)'�F �uU�ʶ����A��3�ťue�
�dnYsx�u}	��Č�$�I�k{�+W�̈�X�e�8��{$j��gp�+�(���4�O �:�x����5�I�?U���jIgf�J7'ӭ���4>S�=���Cx?�E=�9�5��Q�zueT�wOk2;�k(R%?r����0����1MK�;��*A\vPH"�����f+yjD⛛Y��l��#VP�G�cʱ�0���a�3hC�SDP-��1܈f�u��8+G�h��yS!�&�������M猡��?EY�+S��x�pj���
�.pg	�Zr;M����.�w�/d�t���7�R�B_h��3$�q��ϒ��I�T[�(L�Ǎ�5�kt�/[W<.am���8��¦�/�qF��u�te��I�a%���1z@��+B��l�m:Ȧq�)�|8�v§�ϳ�̓�� �jA{��7�c�q�y_�!w^��$��r�X'⪨�;a>���^p���_tߘ�v��N�֘���l;V�����\d���'�K�Z�=�V��R�N� �K>��١"G���z�m7l?Ih�b��A�a�Ô��_�#wU%3��û�N �O^����%e��O�������O� ���.� ����.R�^!�\��� R��5�{�L�Xs������+��1,gs_����ᗤN�E����y���xhz\��]z;q3�_�0Ϲu�d�x��
���^^5���b%���1���X�_�4�K��щ�����W?�� V��/w�a`�����Ӂ� E�d�J 9����g"�����12��e��y����U?�F'%���m%<L�>@ Kxڐ�˴}^P`�t�*�������Ut"`���:Րİ�լtf+V�Á&��[�^�s�X�-��o����CN������_��3Z\�3����~� gɎ�g��Y'8��h����~!C2s�q�?� ����b�iE;�T��<�ca�vBɲ /:���;��.��tWk�IT�q��<]̨�I�=+D�jǞ���s�l��k��o �.c�Vo�\%�6���r�C���ҽ��Ñ��	�炁�������F��W���Ф�xN��kM�h��c���r����0G�.�l��a��a���ae�6�)Q���4׭�e��|��Y�25���[���1��r�rh�%��d��Yný0��N��-�����u����.<�U]�
���o:�%�XS�QK���6!LW��B��- A��U���<��E�O�{���^֡�Zt��4�3���0��Vk��'Yciś�6�T�~՚����aĘXĹ����M��<;�h>F-������<��}�j�@�8�Zl�P(P�ӳ�d�{���⬇��Ѻ�p��:��e�񚍅�N~��7`�CQ���K�I�����Q"VY��õMJC�)Ԯ#b;�e�&�!��d6��=;%f�d7��O0,�˧Q�@�T �a�HU�{��YټRq�a�Z[���FbΉ�r��>BP=1�ǡ8���+��Day�F��1���ѫ�]�e���,�N�N�&XJ���d���w{�Yʝ��F	1)�P_�F��x3�z���qͣ��$c_`���^ b�&�Be5��S}]N��)���L>���>@��Ȭ�*&�
(�?|W�QW�;@�!�Pm1��k���5
���ms�b�^j ��qY1��ljp���B�*]?�.]aiW��bb�QzC�j�_y���M)�{�\q��+�xn� `K�9�'o;����U��d�x�􏐺V�l7�'��K-3��J�׈Ʉ�vA6����~�}��k�}=���l��ձ���r	w0^$��tΓ�h���l����/d5E%�	�&�K�
��]�}�f��g�������M_fX�g�-\sAm��2�D��:hlc�ݧ`��>��˝��U_�����K��H:/�sW�ʇ
����2������gF:~��8��@6b�Yٸ`��,�.����M��V������},4>6�|~��Z�Lޅ�FnKtrK�5ĸ}-֒�.��n�������A��eפ]km�ݪ;z��7�UKה�L?��	���S.{�_���݈P��3X<�9M��ylu��
fQ�幰8���)!�nQ:����C���9n7����uh��@"��~j�U����1�r^7t�]��k�GXsh�4���#��s��6q8g�r��7��5- :_3���B�Q?c5�]�,���VW�����W��V!��N%�l/�S/����쫬jv2�_ؒW�Fl3h��HJ<:6FJ���E �Bp���e�|2�j�3P߆��U �3�ˊ��}_^�q�o@a������!���@�+]g$e@sy��^�.��K� ��^<`�X����n����yʁ�r~^F��#��=�/�̋�WB���P����j������o_��a����U��� �tu�5�%*0���=�����_��;5��a꧇���œ��ha3�NŴok:�}y�Dd�InH!^�w�/�	YԚ�g��!�fy���cq~��[�k9�2�
>I�}��@k�=�9G|S-Y���i�-�Q���%oZ��s�6Ƣޥ����9��ɤd���V�I��v{�Ӆ=ig7�S�w��$�.{װ�7�������@�� *�f�D#�֯��D��R9�V�C�xb��6D����#;��W��Ӽ�a%��������:��"��͞���(����6��ܲ��.w#< ����Z�כ?�=�T�������kq=g�����(9� ���R���U0;N�=t�`���h�E2�E��!%���~*�I*�<�7-�xgd�2J!�j��wC�'�ي?���c�1�����L"���Sfo��f�;LF�9�So�ǉ)�0�m�"G�"��-���pb	l�$���K�",���A7j7q,�\���p� Cj�R��E��JT�}�EO:[��iA�yـ��ZAx�.p���1�V�}�
.^�[�l�}���g�C�oG
l�tc����'�����\[I�;6{��p����ӂ��@�/�xT?�Ao�mN��rEh_4]zD��R�r%�Zdc�/D�I�AC�_��W��e�	��y�a�T���*�j4�@��;�[������{�A���m���%2��OTB�P\���=�cݪO>���7�Ż)��8�)Q��AWA�̛B=��8�J�DXQ���%¥/��t�yf��sh������eD�у�]�����d
�WwX[�bl������Q��i����r4I=9�C6���0�g�`���?Zs60kD-�NYRO�"�����I�<i7���#ڿ�~?%�0�^��2����C�89ئ�� �ѥ���� K9�e��t�R���8�����:>\�v�ZS��|���&���X8�B�,���+���I�J9g�nm�����S�Z�=�3����;a�x���̜h�&��3SX�A�o������%�x/�P�2Wq��Σ�_��(���,��*��I=|�U �tE���JO���u�3�w�D�OM��ղ|����Tt6*�^�$.�-�?|B�U��z����=��}([�|3�z�f�����Im���޳�s��ň��X�ެ�'$9[�o���
0��g?@����^bʀ�)�Q*��8�����H������tr���1�P��>c��ZKIL�X�sէU8��{ĺ���G�U�M������A��Lk��
B�A�4 ��yQ�p�*�7ۨޗgo~��k�2s�JP�4h���p{rnˎ�V��Q�4w	�g�,Ͻ��t�E�N��I�$�.Cȩ о,|���L9��*U)bs�E��[�R�9����J�i$�6^׍sd�r���#|;�p0@�"���dJ.���U�˙��춴/;��K��1W_�ɝ]~>o ��P���wJ���.~�ugR��J�y\sR����`��%�.�i7w�0�}K- +���9�cS��pcG���^�yi��d|t���C�o'�̉G��7�Qnak-��bzAh�J)8boߖuw�r`�y��ȵT��Џ:ak��)���A�K�z���t<�$\�l�^�f�SKƻ ��p�~9�p|(t�L��s��F_��OC���{�|�Ur�ϩ�ZIjĔ��y�)�s�<��ҥ��mVS/Al~>�Q+��G�l:k��2�o�p�:I�y������º�S1�9'Ll��G�pd����`�L�����p�m�x;w6�, C�z(���0R����tkQ̉<��F�gf,Ns�%��|epk%se����ğ�����y�3��m�m{����h4�.#P����[?�W�E6��)��[�Y���
��w٤hFټm�n%����0��)�����<���IZ�+E��a��"��U8��5|H�w��7�x�V�3Xf��ZY� �ġ\�z֔������ ,�iP���}�x	`�-�ѭ��7G�ۗEi��;��t_$u>����wNa��
n	Fk.�������|E%�Tn�P���|g� R�.T<��|1J���Y�����y�wd�xX��v��L8����I.U����}#�� el�*�
�y���d�Y.!ݫ�a

�;�� ��ov>֛y��F���?���p�m�����Z��ٽ'��V��>$��g���O�Y� �p�C�.ͮ�8y����ǹ�[�X���MY�&�;���5J���u07�z#:�"W΢põ�Z�C�����{nĄ[���yE�:=��2K'�/�k�~�3[V|	x�ҵ)����-���%�̕)�\�_�ѥ�����y`+�A��S���/O^���cQ����˸l�,ׁ1��Jt���.k�["ޔ5�40�Z���L�`'"ڹX��jJnɂ���3FUr��W�Pw��J���/�l���q��O���mt���:ߕ�����o�1I��n�@2�3�U!�gPȐ��+����<��:�2��.�81<�j�[?Ԑ��!�3���C9�v�������
�'��� w�L�roG��6�!��=nL�ZD'%� -#�uhEU�F��0!��!o@l�C4�-��������	���7�x��b���>hʅ�v������a"ɹ9wx�wyS��Ybj@`zD�8��q3~�{������jZf|�;���s��r4��N���W�N`aЅdr�v�ε[���G�2� ���'Y̕X����B�`����)�������v�@��! �����&
wI;�8����zg��*���T��/�{�� �e����x�e�Z	�6�/+�j�-Z��F�?�6�S2߾MRBA�.�b!��x��sP
�b�j�C�uXݒ�
ʜ��mraҝ���o��x�'B3���4��=��d��t��z]u:��Z|��keX�8p��aD�BK�w�4K���H�MZU�n��t�r�`�������$)�_��7G���=#f��yL��`<�
j�_C�
�;��������a@�E��$A�� -���uo9�����2�s�{��Ԯji����f�E�ઊKb�_�'ƀe��<��Zb5��ag�ؘ�� �6v�o���\v�6��S�ņu8�?�*����ܰSy�)����_�-�$�a�4�sv]�uZ7G����{L�/lP&�G�����20yN���=]+wd�:&����&�/T�_��C�d�F>�j�/�ks��哘J��"7�8ej��v�wX�>���ū����� F��xΡ�I#��i��V0?li;C�5�1���xAm K�׷� �4h��YW>�Y�����ø2�1�����&�< �1GH%��
P���R�у���"`����{�(�����ct×v���NSɌU��q�t��SG���|����2J-\�~4��r�G���'[/T]�N���%�=G���w�,#/����M����鞢�СΘ�q��&�!�b�}r����Ëtҗ�0�ef��2�fL.N�Ĭ�ݮ7ce�� 8�%D4-̻,`uN1 ��<7z�W��R�v�h��=XWwT�T��ǣ�[]weΗ�N�t�\��R1a�id,�?DX�$ݦ(xTA�4�ЬK�P	��M8@�k�q+њ�I_^u��^x�3=��P��3��,z/���sB;²��c���I0H��;���آ�E}Q$94f�i�)�i7��/��w}�L�fԌ�r%.G�C�<
3,��П�Uo�:���{�|n��MJ�#��x��;�λ>���l��� ي!�| �G4��o~�;�� �0`݋
��,/�5��\й����x�Q~�d3(f��yj`O�_�R���������
�4c�l��w�BdoZ�^��V�s� i��UhGȎ���0�Ă7�y��U����#_�
��x�6f(g`d���y)�3h�M��'~n���U�r�)�`�)�k��� ��N�k@��f��W��+�hNV�c�x��V^ֻ^E@Å��Ы���j�0�����ԾJ�}jH��T�i ; s:�y��1*��UQn�3�ÓS��%r~+A��Ƈ���p���Ԅ��	�5�����%Nk7c�zrAxT�?��͊n��j�aR蔢	�XK�fݲ���XP�)@t�=�&�CZ��}ɍc����u���L��٦ r6��
>��Τ�Q�]l��Ѻ�^���r��k�`@ݧGV`:ǉ`(�"/�7J��d�U�گ���Cr>��+��R��I�ϟf�>��1ù'�!�o
�ҢL�R�Spk�:��ǢT/\0ȌGO��
�$�,���ؓҤQ�6@���`� ���֩�g��cE�s���B4�(�P{YXod
i�P7ɲ�,y���=�.b��[$�J��9[�V�.�2QLU�oP�K� )7��!��Ge潆�k`!�HW�q��V�`�����ɣS��qlA�#"�L{{��/�HBU�#�Ad�kf�tQ�iy���I��灧��5��I�j�?\�1��d��=G��2�cm|ȥ�������G<SX3���v4T��B�"�Ul��^�K%�鼆�NCxK�qyMs^����pi�[���P1�s���}zE4ke�x���c��W��eY6�����ER�=&?���94�B��8����M��R���x��PV�"g��r�e;��Zƒ�~����^���H��W:�Z�[Z,�Ⱦ�i� ��S{^���K���z?`��T�:]|�lۻ�sc�����T���q�IB�iB~H˵�P��k<9]�Ct֮p(s�$+�f����qyJ<tt�}<���c��wU�c���wf��y>�(И?�o��<���D;̦V�~晵R;����0��BxºX�G�_ ��49�ď��^��ٚ����<>�}�Ii��\t��Gv1$"��8T L���X�G/�}������
���;�V|��A�$g�`����� �����)1����Ty�Ō:a}~�4VA)뀾��⫞F���vS�-�+:����.�a������Y"f�z
�>{��4:c�F�p�7��:�$���qTx�EVI��FA� �c��z�֚�"n����Z���K���vm��wߤ6n�4�vE ���xI/���s�J~Ĉe��tk�O�"8����'>��B��Km0T�����3�t��.�71z�4L�h(f����Z ����c�#��C4�h�=�b���N�_*�`$��?��&nE/̠��K8��Qj7�&�,\5�Q��F�~�����h�Cn��4z�;��i=��8��%�NE��>�)��Z#�8�F��x�3_���{T�!���W<����-y�4�(g�`��w����H5T0G�4�P�d�̒h]�`t29t��-->��{�v��߹q��7s���V�G�� )��`hs�s�ǡ���Ք��޴jp���5$�� 	� ���������o>�5ғ���v�C������k;��U�7`��PN���&K�-}(/���N��C� ;�;�[3|������,Z�I�t�u ���E��;��+OSM�`^-nmT�5I���Re���d��FB'�����P��/Ex�\�}=�_�qBOJ�́��w������k��$kZC�_�0�T�kyX�B��ܷ��h����~�_�3F��I̹�'��|t�?���q��!u�����I�%Y���� (��b ��݉��El�،���~i��z�ZP\n�Y��Xf��砚��p������?�	���;��>Z.:	Q��UՌ���\�듐��t9Fc�e�4����r�_����خ�#X����w[���qz�
 ���H��#(k�Q��0��e���� D0�T�\�g�c�D�X�����u=^�	�a1a(5���#Y�$�/�պw���f/�*�ǹđo�r�2���"�&h��#x��G[-���D��Q���%���zQì�fA������/�\���ʃ���`�����K�d0B��Nbz���蘷2(�3t����X�a���Ϡ(	/������۹qd�<Pk��}*zJ��^f.�|f{}.����J#}��C�bO�Ց�م�C��2S3���ޥ���ZJ �n?ì�cL�ǽҵ3��9t��\`	�^��3�'�;h%vou�j�!V�и��#J0i�-��������ѻ����Է�pIo�ԿO:<)�bǵevy{`B�n�\2׎��zi�#�G��U�����H�,�4�"�K^��@j|��
#� �¦)f� �h[2�Vb���]�=r�f)�w�h�+���PH��2~n���s:n/�qt�.f���B�)l�Ҡ�N�F'�{'�I��v*��T$8��?�GDQ��24�+Fǰ���4ʉ+GdU��%g�!#=҅�`���n�b��TX���]K�bK+�J��OO�]�l-�(� �ҥY���g�Ѓ���az� >�b%Z1e�l�♚���ɽ?��Lwh�~탸[����"��%I����(�cR�0�`O�l��;���1�ym�H��b4���3�[7@�[�XR	�O.oKs	�6��.�z|AwF��݀ҫҨ�R��e�y���%|�O�Cm6���>,�ҕK~�=Ռ7��*Č@��/�U�<��c��՞[��nդ����*4�'�e�hߧ�o�㴽������!���uЅn��jC5[g'�t8�pƿ�$H ��8;�(r�����c7B,�9_���(C`mƱ�,� ���aٴ�f���3A�?��
1�D����Eo��9b��'}��7^��(?�Ŏ���c�,�E~���[ׄ��Y^�6���g20�Д]cY�r���x�dţh���{4�(4}xN/�k�5�z���{����tS�h0�A�XX���{�A��ar܉�/��N�~�}0�{q�c���=W�w�5JW6"���Вn�j"{38�A��d�j�����v 5�͸f����i�H����F5u�KVâ6>J���@(a�!�B�:�l�.��k4욶��.��.����3
=�h�"�S��#�� ��.��%�����D������"�8��E��}KZb�U���tX4��O��Dޫ% ���*�7�s#dN��DZ��42�,��FW��^�=�?����"��xS���)/H�+.�U��=��)�� ���z6D!z�?D;6GS�|�w.!_�ړW������g��c䒍U>n%�fI�X�{���f�s���UDʬ�Hg�<�z\IU�M�R���nӝ�=2S�&s�Ǝ�֬�@U�:I�귗R^D$Q�ɞ-�l�93��n��;���K[�Z:������Űp�<�,F~ݭPL<�p` ^�H\>sS�;KW����k�t �X���@�Ǘ^$4��Պ�W�Kkr�P���v�����u�qm����Z��\�h�����o��9nV�u#Ed��T���;�0o�_��^߿���x���׸/�	�Q������RQ��|e���9���ZcNu���T�tWǎ�Lj+q�A�����.LO$��5wJ�B�����$��le2��}��&��v	Sd7Ӆ7����?�_����ZqT��H����|l��r��$*�8��ho��%+r���XR������F.�\O��;�A��w��-���u�⧝�Pp���+��a��Mr����w�ZN��2�:��[:J����?���/|~�wXׅ�F'�ov�T�h=�B"E����g��*��n:��.�b)x�.Ef����Jn��32�_��-ݺ=�ޓ���=�����5 ��+TG%�� _7iا񾜉ӥ߇w?��K:���6�G�,���@xf�`,|s�ګ�z��m�F�3@����/��1����@LJ��
^f�'�w���@��5S�޳��ρoZ+�]��ޡ,�wC~^���O1rd��]�S�����1������1�z�(�Bf��^����ebl�}�I��Wz>h��kG���{#�V^��)�pğ?�	�F3�]�q� ���n/��_�_����S2L��q�!��s� "Qn2P�~�Z�G��U7�5���⫪)-����?���i�F�]��#��^(ē?�����|`V?鵿\��t����br��`�r@�����.������!j�~�qa#Q�nl6)3Bqp�1�Lh�t =ݒWW���\����������($=�q�O�vq#�+,�,1v*�y�1ˋl���औN�ӽ�����(CAmLf�)����5!{�Hז�����د�rW-��.����<��G�ڰz�.*Q��6��&���G����c��>O��a���hi���K�믊>.��;�;�U�FSO�X�Bei�bY@��K��/D����ߵ���O���$W5^��*O�B�3�z���R
����ލ	շ~|���;7_�[*���k�Q���!��ۑ���̛�"R7U(F��
���-����y�vτ%�ߐg��X[��������l�~��)+��ڿ�W�y ]s����h����7�5L�\5�BC��G�(1�i �
¢��Z�z�5��y�D\*.Oȋ���.�?���J؝:^��)PI��U�?����!.L���E�K+��g"ȣ��3�i�J	����-PH'۾ïM%J�� �j,���p �>��H��/g��i�:Y��z뇚��ֵ��aU���e�eo+���`��8}7��qS��� �G-O����RF�G�k���2յ�TE�����d��r|D�W�SY���P[s�
��}�*U�fCԢϬ�W��Ilr�J��0X��/&^>+i�v�qz�]hMR�k���q�����C+KL�8E:����w=�o�|� �"�\8���/�(�8�� j���K��X���5�j&�rt5��p�x�W��ȨZs��v�=H���)C�c%]01��3
�e�6Ԑ�E�%�����m��k�d�����n��V�Y�&�xҢ&t��5�!�B��[��t�>K I����f.����X�SE��E �q���q�%M��#2�}ٍB��آa���V��9���|�j�[����^g���/��v�	���"��&��I�ߜf���P��������}D'wc� ���+�ʰ������ ��J;=?�YP�!Pr[�����mM3�P6P�?�&
B���=���J�#�"V̖2b������}	��a)�Us�7��F<~|[��_��V,�gwut� �t3k�~%(��$�3|�)�KV1�D�4���Z�T��R��1T�jT�區�����}m���[_����Q�W'>�'�'넱8�2拟e��_NF�ȧ��1b�eK���D�����ԁ	�.�%�kM+	�՚4�;8�i6Sջ;e�����#��+@�D3�oނam`1�/�"~X��d�푼�6b�F�c�WX����F^������qQ��3�]+h�����l����SW��6U�����3
�J09%�����c� {:�`<()������I�C�E�'�F�\aA���SV���������E�&�����9�tnߋ��C$��D!�ÿ�1���Y �6GW��G�������ߘ)�g-y[�\�z2g([L� �]���P��i�4|��0�����u���`��A,ɗ�l�jlh����Zo��i���M�����Gx��l�^��׽����Frz�:%�1�˗�Uj�d�� ���^h3�m5έ�Pt��A׬��Yc�����ɣ�Z?��ɝ�;�_b 5҇NF��8�E>Ή�#\�k�:aԠ1r%ۣ�ޫ���0�/�ܞ_%��^oݓ�Пo�
͇Ցe�P�}%a%ӗD��@ШW��Bwv7!��.�&�r�'�H,����]:M	���RI�篐=��¦B&�Z�����U�Q*�U�x��ĭ�0&��3x-L֠�K(�UE3�#����/�T{�_�ݬ�*#n�>����\����U�Z@�ԓ���-b���A�#B�U�]%P�S}� ��u�=�dbg�ぃ�slF����t[-�J��a:b����fM=@hcRv�A7}�u G�8nG��g�_���mQ���mY��"�k�h�C��왕8�˻=-��e�&�o���#���>+��f�� 3�3�gдo�O�k��1	͋��7������K`[(M����_.�uvv}:�{�|�27�d�7}�����o�~Nً?k*l�Ѻ,	�{�:ky�����#'�z�B��c��ƾ�,��R��Q7�6_��E������Xp&e�C�)a���35�x+m�u�)�4MJ���ij��6�ج�^P3A����N��6bx�r2��w���n�i2v�b�ŷ�-�t�n�3 �/@���݅��AZ�Dی�Ι�E�R���D���W���/u=k�Bp�D���.�J=q\��tt	�qu���w��I�S�R̨W���e�%��K_�OH�,��I�#�"U�`n~��2:||��*|Xq!Y<��]�B��V7\���'�3Ң����4���S���s=��0Z/	O��p �Fz���h-F6
|R��g�K�9[������6�ݼ��"�/���q�T�)2�`M�VE�A�eD���UʮY9 f�w�O����H�[m0i4[)TQ���$��H)[�����QS|�i~�!�_�k 3.С�e�9c-�`���+�O�X�Kau�X2�+}	D�qDt��n�?@�� !��bTV^��l$q�Aú9�����E��V)A֫^G��Y{s�X2�9v�2#����'�GE�OliR���A/U0����56F.�$��
�>qA��1P��s�~rHލ@WE�W�
�:٩ؙ�&/�ʸ��M.9e�sNN�vǦ\�*JT"7��IC���G�^Kſ�1;�8.���2Y-#3YZ��c��S�Y�r�xˉ�~�zlaԬ[�^տ����l��iJ�n=�n��0���tkڒj_��N�|#��m� Ђ����Y��ܦ�'{��r�~�����s�!�!vX�[8�"�תu�q�d�q����f2̳����,u�l��<\�V��g~�9A�Dv�L����U�ko���?1��4��[;M���^(���������Q�gE�:N
^=�����]�uQ��W4��MV�TPX�f�$'P�f����� '�ά,k3�E���E��N�b.�	��[��Cv���Z'��|��K6�a�-�r]\��Q=uOKd�[�����ʔ@������q��ȣb��}�����y!�K<�w��+�<�"w�ʢq�v�mq�0P|Q]�Km ؄�g�z�e�Y��[�<K�S�n�[j�ј�^�-q�&�ϥ4��4ŧ{�X;���˞�A��������0�����J����j��~d~����ZwN<�Kp������'��ð+eS��y��Obn�Pː�h�p�.�՘^c{�]H�Cʔf'j0Lp��%��nh�2�@�OC쌘�Ĵ����W�lڗE�J�&�:8۞M��	~u$3���?@���2|w�����N��ߝ��o��'%b�1����=����W �Yb(Iy�{B��ÛU��E[�i��KA^(��2� ֈ����İ���u�����o��Ku;�<f����g\��Z�)Y���J&Ƥ�hB'���xN��^H��1į_$L*�iB٬F�m5:L�����2Q����'�f��C��ozʪ]�7�{�� q;:�\/L�� �B0B�8��.M����}�Mn�M0��@a ��-N��Il��C
x>sLm	r�5�W >��;9�r�b��ݒ�TX5��Y��}�C���Q�q��� ��Բ�7�f	��K���C�/P���!UT��1��
�#"5�0�����c���ۑ�a6���;����0����A��u�~ư��3�M�B��.^��k ,�b�Az1z��R��ÿj�����eu�|r�b�L�6�����8	4����%'p�����۳n�)�M�ܶY�Y�����9��7X��뢓�,wÍl��XsR�9�'�n�QH���kkJ�|�G�]�Ȼ>���9��}�@L1'�%E��14 ��ʟ���9����&�����@v0BK��(F��������{b.~�0qD|��tb��"���B�Kʷq������3|-p�컼[���_ښt��;���aV/a�a�ޏa=��T!�d�N�(�\�!Y������Ѕ+�v��q{��jzU�j��I�������	v^8����}�c�I���V����\bAmUr�����!�������ώ*�?�a����1����1��3F}1�>0���Gn���{���~�{��(�������n֥�>(U�Ft�?��@�DPm��sn����ݝ�e�	v�� t�(2AKD���<(5�X��`Q��ʧ	�=i�7]H{�Ѣ���D:=��(V���ɚ�I3c�+��y���$R�	8��q�Э[9HD���s�Yq&�WPF��%�~�%x�ݞ���mW�%�D�`�
Q~pg���U���� ��e^2�543�)}E�!G]�#m�K���J|Ç����p7�~!<z*�ƾ���\�4e6>^�����.Y|���>|K�W���u�0ū���,WĚt<���ɒ�a�kඤ�ͤ�r���~h��;[��C��� %6t��3]Վ#�k�v���n�s�|��6RU5��W��d�Τ;���ח��`nDЭ.@�>4��R��>�T��t�3��j�-כyI�_.X�C�i�}�A5?bd�Bb9p���8�`qE&$)��E��}a���m����*o�<y��6`��#WGR$i��O��1��x�'4n��'m�6b��ۮ6�A��da���H��Q�c�
z��x� r�n�h�6_?�w�� Uf�=���įU�ɭ[P��(Tlb��`��<��6�9��g�u����b����k��_E���V�N����X�nI���n�M��[��&��f���N��0[�5��l���G�]J�(c>=���e��^����ĸ���>�`H�鬨��2�����K���o1tڃ�=��-; �qp�����.?�=�ؾV�����o��A�k��$&N��k�[4J���C_�����f���7I��~PC�Σrs���3�`���b��Ņ#�����MqB�s���p.��A=@tG��S��Y���
˕��&C�[�H�ڀc]�L��b�ҥ
3��g�R.v��u&OϟPs��gq����z��.�������+��OpR�4���A6�����Ӑ�e�%/$PS��[����-�HVd��b9t�uܴ��H�:L���k�������|���S�+>���Z�M�C
�P�L��qHR��y�Ĺ(���#�t{?�T�����؛$�����3�1�QY�"@����@1�Ƹ���B;p0㋃��:�����G{}��(4z�.m�(��j�"��$�l1��1��rh�3��J�$7�u�f3��
t#b��57��;@�r�rҟf�W���A��ظݛ��i�;�c���b�g���@�b�!oRKF��2��7
�E�ėXif<Y��ge|.A=7�dg+4�
��zh ��u$�����%���3иh��@���λ�S����P�a�vu/u���L��z�����2���Z\����w!�cbYq�_� p�����S�(��J��K'�l��·���f����iײ�C/#A$�Ư8��Y�8�M)_"T2W՞k�al�p��
F� ߚB��q�M�B��᝹(r5$6vvZ[�Ś(�5���NZ!C�?Es����B�y:��gg��0�K3u�i�5��;�����YׯH�-�����:�:�M ��y�n�OJ��Q��~ÙE�2)/iyR�ġA������7YfF@�����V���<7@������J[;}*����������";����Kh�r/І`�%+n�\�����C��Vv��w]�7�F��?�N(��n.!�-�ѐ� b��A.G�9֬��Ȇ�[�x"w�3Z � I��\��t�t&��4��~@�«)u��,ٷR��� e�O?�,�Dv[�Ն��1~�H�Ʌ�AQ�k׭n>Q?�>��G�d���]�bJE
�ر�h�2��'�0�76���X$����h�ڐw������t\���b��y�XO��K�ܢ��̻'�
@o��W@�璘��z���[�*>/z~�ó�q��D�!�Z 7u�s��&o��oZvoD�5�2uO�͐%	Ǘ�^ϐ���=_+f a}�|�'@mAZ Z�{k�{6�~������V�U�]��_������!u;'�[�U������f�_���B���{�q�yW���E�B�-��M{F(�b-�>{���ѱJk!/����S�\�M�)8���BET����{ѸBӧ ���3mѾY;�n��K�����V��/mb�p.�Kc�=`u����S?(�O#�L�̓���r��u�l�X.N�RnD�	}��ky��.���ɴ�ଲU���!�X�����-�ӏ�.�,��3і���2oDv��z阫j�4[^�PФ��^e
��ӵؿ.�t*���|ݠ���,�|f�W�:�Ё+ۼ�9olF:�捀ްQ�%M��(������#�K���/��,	y����p��E�Aj �^F�Y�)A�l��mu��&�c�g�Ђ!���܁��|)m0�p��/A4d�bϴ%�w��(����^�iV�6�i�w�Sc����Lhz�g!�R��I��$6�����L�4�">��+ �HL�D�ER���Q��i@��Lބ}]�n�- ��bB�fN5��lN�$ϗ~.��ك��B˞Օ������^��CP���p������͗�T��+;L\����Xl���m9���~�o�_�C�*^*�0�ɥ�
�0��.d)�H�ص�i�����k]%�M�������d+��$���e��;s�˪OH«6o#��Y��*���ɲ&��mg�(��<wy,��m�%1��Q_����%BD1��Y!�k��eų
�h�@Z�5���ր�_�*nfqF��H���yȯ����i#}MR��UjY����o�����|�Wi�#��|��ߵ�h���;�4���I�Z�(:Ö��Ts� ��SX���JZ�S���$���v�\��,=���׫���e�j/�����Gr/)1�6TvH���ČE�Uo5q�a�H�!YA%V������e�Ÿ�[ RF�^)����������r�Lu��=�EE�/�&{�_8��E�����a�L{L��V�Kv1�A[��@�hw"��ѧ0(vO
�[�q�X�2�Z�6��e���G.@54 ��߻e��"��	�LYz&WC��^s���>�;����+I���Q��`E)�����k�}�c�c+NP�v���`V���8��'����h(c��{��7�[t�L�3�B�-&�@-��M1���@cb�D�s����9p�>�;�;�|#K��M�%���ɦ�V�gEq��+�\R�O�Ͳ�׻'��z|��D�]J�̓��Auf�'4���[ߞ����w�gԆ�~��YQ]���G%nTǭHy�V<^�p�|�=Ԙ:�L�r�>^�b�R32P���x��|7N���
@&ȜW5G(�u�Q��E���#� �ޓ�ib:>�I4����9�]Խ��;�0�݊)�Y�_q������K�����O0���uyS�벤GX ���c"�B�2M�9��/Q��j6�)��?���+Lg|��������$#$0�������2Z�I����K3ǻ�	W��� ��}�CwBEZ�#=�]���(̮��r;�*������K�\�fV������YT�P��.�1$���.�ߝ������h!R#��v��9�BP\���;#U6
$S{O���C�)�2�"�-��)�{���I?ܞ*�4�P>��h�x��U�yo[l� d��]�In �I�Qcn2a��v&�C<W�ί��~gm{ Rۛ��r�ƭþ�;�$��]m�������� I����3��jsJ�~mM*1�՜Ƒ_�B��<�����=)R����ݫ�LD�g���;���= �:	s�N���kt�?&��&�;W_.��(���A�Q���02�rc[��	,����1���� $�ǥ�ʴp�.�S!�!A�@!%��gg*�ȼX=��Az�ǾE��&��VM�B��3Ԇ��2��5p��X�}���B�S	�u�@�ҍ�;����5�ʛ������,���|�u��8�"0`p�L\��� ���vQiQ�6�@u��V*� ��huU��߷ެZ�8���"��n�!��%g����U$����5Ώ�I_A�Km�-�{[�ޜfT�pI>�L.���n1+��J��9����ڒ�
�U�{����$� -�!��"I����C��d ����T���&����~+�R�b'QxW�e�w2��\
9
7<��Bj�" Lc��U��"���8,';o�����s9�`���4�c��9�opVB�Cd�E�JQ`�"W���Q8r���h��uWv������'o�ux����h����5�WH�dZ����̏� @]��ױ	(�2�a�O0|�264�#�4"�n�ъ�~%��h��b"4>����K��Kf���+��.����bDr���pc�?���h��8ºAuo�
I�r?�+�������؞iY�������>0�$�
Ͳw�t�p.c��K������[~��kB���P����7jE��|�����޺��ˁČ�n��n���V(���~�)7��@4��-s5E���?��n�ͤ�Kg4����m���%�Z6�b��m��%gve���bO����g�*�]/s�{f�Hy�ǹ1p���R�d��[�c�
�����8w ����1��F�?~gg��,�n�(��%�5B��`Gq@_#�".c=��KL�aFƅ/�&��:TnA�c��\�=6$�JU�f�e�!�gY.�|5XN�Oc�\��#�;m>�Va\8�u��ge����V���Fz�u}L,/��Z��e	�?!��HӻGs<�z�5=bx��@�րtkTY����6O����I�D�r��i���B�1�}���c�ۇm�~Ȋ\E�#�n���5�����_��_W!�B�8�lK���c��Ɩ�i��<�g�A��2&Q.��0�V�IE�0��G|�_�؄���_�2�TO`�b x�����@P%��L��������e
��c}s+!,���e[�N����v�G�0�7��k0|3���\�ͣ!q�wyD�X`�β�щ���~�}Ԯ��
�x@��[�J��[v�6j�R�Uˤ�?���ۮ�r%��!�%��Ѳ��E78h��ˈ�tZ�r��Op{��+���>�\�'�
���؛�c!������0>�F)57$I���Ra��c� Z�
$�A�%������඾F�t[Kz�{�#ldɺΕ�"5,�^�k�p��2&�w��lo�~��$�b��.hjD&�L����+s�?�J�w�{,i���q���:����H���I�0�td�84��.e<�Li+��B�Bq�"�q��#m*��E A�G��g$��$���P�^~�|<ŵҒ/�s�=g�g1Ҝ�ͼ��Ь��Exc˱ev�����+y��n0ߧsA٤w��>[��u���g�C�ד�:k�cҀ��w����6#ɽ!	/�b@�������%X��E�[䵼�wH�>�J��6J�%��D��c0�)U{�6�LC�o7�t~�`�) �O�u��!ss�!�\�v��6cֽ�>�9�~D0����Z��D��c���b�^��~:>@kI���f߫�F�W�'�.�bM�%]9ݗwy�eM��{�W����7LQkM-w����Gj��+a��
��� E�L��)���sЕ��'��ZP��I�,��-��G���H�Q��?����Wi3H��P�P���4��Ҫr��ˊ�T�:�^����>XV��r~�i��_=b΢A)�V�5X����M=t׭�o�6`� ��֎��Dͅ6��q�Q�N�.3�i��p�������;�v�/k�����5{ٿpH��>�B# @^��A��D9�>��!�B?�B�U⒫��|6e��
�Z�.�BJ���c�ţ�\�T���M����u �8���y��������b�-d}LP������W�-�?Wxi����r��5T�����C��tyG�؄j&�̢?�e�	Z�̺��Z��/�����!z"��Kx����g7���*�rʲ�+���<K�n�F����*���p��3jN�[Kq�a[�������c��.9�D��GC>��_+�2u���vMY�j�? �+Y�VP��ּP�߽0ޑbHLJ��	[�w%�H3y�k����$s�U�H�#oc�G��L�7��Gq��n+Ć��#~��(#�3p�[�JZ��ˁuY�f�܇�4fB�o�hB�Z��u�B�<����J5�!��0H�$w|�15c��(�	\�5=��rd�	�P�Jó����1t1���`�Cg��Z�t�oV��b	��k�_]FH�wx*}@
ݦV0�t{ޘ�.���x��ǚ:u@�,��h&7,��S&bc674�<��1<��DO��f,�ܭ�g���_,�|�=+��W4�$���@g֊xP�����,��K����6��C t� ��Š*v�NJ-m�+��M��6�HI�8���P��@g��N���?���q�b�X3��q�	s��H��!&W��������9C?4�"����+��8�7m5�O?X}�՞�B�H�p��7�O�^���"')tr�S���׭��&SsT��~&K�F�of-oE����� ��G�,A�ik7^��5x��}��!�N��R-)��/K�m�kd[�j��e�8�*����XO@QhO�A���P��eX6�1��a�Յ�Y)�*�� [@��K� 5�z