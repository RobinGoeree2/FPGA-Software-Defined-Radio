��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���G�H�ƻ	�"�iQ�����3�7Q��㼫F|�ݽ0��@h ���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�[@�qR�� �����t�  ",�N<��;���Z��4d��{�
��|��Ȋ)zo1���á�rezxB���]Zb@�q�*�+
MہW��K�F��1�:�Ω�[@�qR�� �����t�  ",�N<��;��� B]�pE���	x]̃Dj#^Da����M���Af\O��x^Q\7�z����)�,�˛D��w���旴4�����<��a��rl�ʩ{�Bf��� ��|4�VDG+�������X".��>��'��E����FȬ��"|���2Ee�Y�R2
�I.��	���
�ƭ�IR.ux'V�vЊ�[-c��lJ��p�E38���E���2O��'HY-��Yk"1/�7G��D�:`�'ࢯ��(�R4�K��9�ĒTC��0��0�\[Y���c.$��@�I��c���Կ���PГ����"��N�� <9[�8@������G�٘���ty.hSN�����\�4�sP&�O�S��2S[����]��wG��D~ƅ�ߓ�7C��H���0s:?8�+4ԡFZ�p�)�3�:_�r,6��L1��m�!=�y����h�},4/�0��ǧ`ZO:K����c�xi��u���;���!r(�J���^F='���cu� ��o��3Ai7����$�c���A����������RL�a)H��dd�@=�~篟|�K��l���y�W��p�8�:r&@����:8E���x'rg����4@-�`\G��.��W: xt%p8>.VVmCu��w)�S��X3�� 6��.77�ƔGІ;���{'�J�Й�m�@�5� Y]�ߏ��P�umSe��S�7�׫X@SY��7��c�y�![�$z7��+T�Jfu�Z��"R8�������ì���Tl�
� �AH����Z�~?�(�Y���m�W}$�b�k��n�L�����Y�b�Cj�,\ަ�It��vȯq�
� �AH���2\��������U�7��W/�HeБ��X�6�~�MUs �.Eٓ�9�:�T��|��=o����"���	x]��:Qt��t2Ϣ
[FH��C�mbg��x�T�o@���q�&E����}@#��"�Eiu��w)�S��X3��¸��|Hj`ѻB�/o����qE�J�Й�m�9�l�U��ͦ��^��9�V��r������=�kM4v/N<E�����C^�Lc�VR���"v�D��"�Y�
� �AH���н��Zk ��U����GW��zQ��n�~�MUs �>�u��8�����
���ĺgq?��ᨾ�>B�y�5A31����(����m�!=�y����h�}`29�$zFs����h5�2�	��u���;�'�� +�ۛ���p<�������,�\	ڣ��G��st�(W������R��c^����s�}�(7U�
� �AH��KH��Zk ��U��:���R<�*:>�~�MUs ��=�����r�!]kg
����?�m����� �x�"�$�Z�G�:y��t�jPP�
� �AH��%�i�6�KZk ��U�i��-a�s���y҅�~�MUs ˙=�=���f���e(�܀Q�ӎ'�d0�(""J7�1��%��.-4����] '�bJ�~C�an��N0r�O��C��0����bm���?d�!*r�/?B�myӖ8O �L#6{�I"_�wms,��;�Ӏ�AV�R��:ۭO����Ĉ���rl�0�(�!��#U�DN���IR�?J��p�E c��(�U����	x]̍�9��HB�1Զ��B���b�C���)�$�ɀ�&}Xa���������X��(��n�T\�G@�{M���E���k�8���҆�|n���6��.7oP�[쐍C40��w��J�Й�m����
|H?���v��EȈv����i�	�����;�u�2�"�/��p����RP��̰]`��*����	8O�_��u��RL�a)'r�Ӟh� ���G�/9$�ڐwP�����Â=�7C��H!��"�Y¶��1�0B(�� ��ͣX`��_/�5����`K
+6��R��l���1Xm�!=�y����h�}[q���%g�Ǳ���N��D���fo?�M��;]�`�}��_����Qr�O��C��0��`�R&.1�|(G֓�`����u���;�'�� +���9gX.Q�3��<�ؒH�ԯ��`�bq�M�40�W�wƼ�=e՝���bm�!=�y����h�}��<]~8+|k8ZR������w�0��o?�M��;]��Z�F�ܿt-)���T_�i(넃���ٳ1P�f���g1S����AX�0���U�r�N�Þ���k�8���҆�|n����e��m*�;r|@�b�؃��em�J�Й�m��JNu���]�ߏ��P�umSe��S�2�:,�nr#�9l$�/P��pO�c�c�ENk�lAc>b�G��8̀@��k.�"SӠ�|&��c���m�Rܙ#l�%q�M�4�}�����r�N�Þ��t�U�PD@��k.͇�@�L�v���0�Rc=���T�1�\�^6uk��~1f��t�jPP�
� �AH�}��� ���'�Wا[��׹�ܤ�b7�|�ÝF@�4%�0�iN�
_���*����	�U�����0��K��l��fu�Z��"R��)F���b��\�4�s��{��]Qǯ������k�y�-KS�#�(9u��~�MUs �>�u��8R���\D�	/E�CԵ�_�!���<< �sN۪�c�	u�~Rp�,k���%k�&ָ��sE��D�őⴔIꈸV�MT7xB2I�d�HnULkIh��:h
�[ϸ��W�A��S;CM���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcN%ڤ L�y#��=�V�k/c�X5$����ڼ���Âﯣ1�o��o����J)�j�n@��	��꦳�FZ�X/*���U�݂�ik2)�
}wʭU&H�1��8�h7H�u�ÍeRuw�C?3d,f$�7Q0�"<�F�ٴB�I�SbW�{b�2"���Bpш�#w��s8[Z�xZq��t�1�:�Ω�`<4}��o�r� ��J��ݪ��Ny5��	g�y�+��T��C�NJ���1�:�Ω����	8���/P�p�<(�P[H�������'SR����.�}|��ι%9T��7���S5H�j.F�6�Z��'i�tw:g+��T��٤�2[51g.� -��E�I�?g�f�$��P�`
5��*�z��Yk"1/���qH���Ny5��	g�y�+��T��٤�2[51g���i��T!ea�8���*���g S��/P�pݒW*g;X~09h�i�k1i�f1?�e�Bw�M�?_W�\I���A#|��[�m���w��L�����'�@���,������0�ea�8���
ae���K�������U�̺��t�iZ]XF��������3bQ=�3�� �֤D�A"�,�>E���#�ڊ<?@��[	J��;��2�F�P&l������g����=�Q�^�y�zL͊�q���{����w¹��<d���<
DN�!�`�(i3JHn��z�_c)���8�+�p}>&�&i������ ���3�ҺIÙ=�H<z,Ҽ&�jV�{+��]n��!�`�(i3JHn��z�:3�>�<5��Q�[TّD ����R�^Ƒ�� ���3�ҺIÙ=�HF���m¡�L�溥����v�8:.��w���\�v���GAџV��0O���ġ��,�����l0��F��j0�T��:��2�F�PY~�y�����[��Q�^�y�zL͊�q��UG�s�����M���HaU$kX���g����=JHn��z���G7����Q@��j0��yb5������i�%Ah�%4
>��XP���i-�9c�,����<�R_#��-?��E����F�Z�>)�����˟y�t���\�W+�[Z��!�`�(i37�ܥ��2����*����i��>�`�0����%����Q��K�����7�ܥ��2����*����i��>�`ب��~��C�8�J�Q�������i�7�ܥ��2���5jy�U�5CS�|i�8֩]=$���Y��)�.����JHn��z���G7����Q��6�A�C�r�X������4];ˍH��G�S�w�Qٶxp-��wH�HͶ�i)J]ڟߍ����7�ܥ��2��x�ǣ�Ò�ÝZ�� n|��_x[>&KӔ�o�J���" (�P@L0��U�b9���:&�>��sN-Y&yo�q�A�o��d����O�]�!�`�(i3±�sR�{F;�f��X��Ye�?���j�g��$Piq�VD�Lg�q��Dv;gJHn��z��r9�3���(�ʉ�I�,B�����B�[7�d|���XP����G�u����U���g�թD�[*q"�?�G����8�TP�T�K"
���d�8���obzĀY�ɡH�� �YߥթD�[*q"�?�G����8�TP�T�K"
�Q�͹�Ɩ,���#>c�0�وݰ0|]<w:�"�,�>E��4];ˍH�F�n�ܱ�7̧�����A�����y������i�!�`�(i37�ܥ��2��
[���p�� +@���a
��|���\G�Y����-�,��Lt�2�tN�By3��<�]�!����M[��Ǣk/�z�xEQ�����5	���]���>����C���"����Y%T��BPe.��xu	�>��l%i�-\1��pz��S⏸[��c��Et�Y�{'%s�h�v���5���T�`�|��K�z�L;Л��Z�n��[��{_8�Y��=�}�Vݨ��������P���Qi�]2�y�Z鎬�����,�q�����CsYl���#�]�!����M[��Ǣr�x�e�X�����5	���]���c�A�L'��!�a��5�%]���a(􆿳����^��$���]׽������E��@IE�U����S8����;(���5�%]���a(􆿳����^���#}�{�,�k,^+a�@IE�U����S8��$FW �9�װ?�p���5�%]���a(􆿳�ؖ��d�I�� �:&��I�?g�f��m����bi�ī*����1�Wa�b����y�E�nwE��S��}|��XH�����,>$+W��� j�(����5�%���(�-X�Ç�eR;�{m�Bk������h%��b���ò���:'�>����߰r�~;�,�ތ�@���[�Bf�^:�8Ϥe��b9����V(�-�ǈ�A0
��T�B���3���ne��'�{�a����'3:{%:k�a�2N��n���?���^�ތ�@���[�Bf�^:{lGD�V�B�M���C�n=ٟ��@$��6�[id=��¾ȼ��#�a�Ą�`����z�.V���)�P.��� h�ҩ��i7N�_�#�6���9G 64ظ�ǈ�A0
����m���Yk��౉+�+���_�R�G����l��q@C�x�>���� �P��#��s}������!�`�(i3ܩ�9�d$��EN�����.V��cd;�K�*A&-�Ri!�`�(i3��1���h�"��
���G&6�+9f�	P2;d�l����O	a(�عH\'
�:qEpCt�w#��@�bR�Rs!�`�(i3�ݚ�Н����F��O��;b�-�2�Ct�w#��@�����$f��_Ub�G��VO�����3�}@��9�ڮWbAg�
d�m-ܐl�}�1�26��oQ$n�ti��|�@T�^��/�/m�d�ů��z��_#Ԡ�����\�JHn��z�c�����<�W�C%���6V���~�26��\�o�mW���'n�^0o�O�A��~������Ƀ�.��|ȃ��q@C�x�>���� �P��#��s}�������H������R\�c��-����f���Ն<i�LE� R��uL-���N���kb�r!�`�(i3ܼp���dkF�+Bd�[ߊ���V���!�`�(i3Ƹv��*Qx�X�ݯ��:5A��pfĉ>99��A0ok��fĉ>99��R�Q���~��p����$f��_Ub��7��G_��'{w#/ B$ Hl�]����g���$6>��m��}�	76�&�j���GpR�@�6�֐����o���\�s���F��������開�u)�L����R৘@��a�\�������޳[��g6�w�9\S�HE���èV��a��� ;��R�ʞ�啅E�@�;���XVN�Ϋ8��K1P���n�)�𣈈�zNc5��;�P�t�5��q&����$n�]g�$��"��є�'��A�:QT��3��Y��?	/~�uJ&��'�B��:ޚkgT:E�DlD�u��bP�9���
��\�v�.$��$?sT���u�I ��d�k��m9{��}�+�r1D��y��-ڨ M;v�u��j�_���ˑDBD���{��fn����3���ne66�v��G���V>�R<�2N��n���?���^��b9���:&�>��s��n4s1ՃV5+��:�M{��������5����ߩ���I_�(�Դ)Q?M8�f2$ Hl�]��Tx4T}����(����W0�]��x@�������a�"�_���3�&c`s��Q����Rn�pPip<ɯ�nv��2������開���Y����Ů�;	�nw(��=����$?���*{ٝ�,���8! ,��e�ŷ֗�e�a�i���S=GϦ-���+���ߦ ���Ǜ��4y�ӓ������ �V��x_ߓ���>�]�\�v�w�?�b�>��}�+�r1D��y��`UNP� ��b�FP&���x�Źx��4�o�rޡ����u>�|�w�佌�&��/Q�����Ƀd�#��Ӏ�`,9�H�Wu�����Rsb�d"L͆�#<W����Yk�����6�{�Pe�E"�I�;�q�hz�:pF��w�ݚ�Н���1���h����˟y�	��x��ݚ�Н�����*%�d�cA�_�Gn$֪���P����p��ݚ�Н��<�I��y�f7$=�0*!�`�(i31���~����l��M�r!�B/(Q�kŕ��QH�RtV�^�y��j��kj�����N�
\�n/S-^F��]�לԣ�2Mx�m�ڨ�hծ!�`�(i31���~!�`�(i3��1���h�"��
�9*�����
�:qEp�;�P�t�5
�:qEp��sp��xF�mJ�0�6�fĉ>99��A0ok�?�JY�)�֬w�J%�H���3�}@��9�ڮW�x_ߓ��6~ Q���L��O��݄�$��F�Ճ����n�~8���a~�d��"J�A��S+e ���p�I��'�{��Ń��Dt�G_$�n�>߻��]H#
ZM��2 �єV��߼
�dgn�*�Q3#*�ۍc(y9}LY�\66�v��G���V>�R<�2N��n���?���^��b9����pP�o���n4s1�h�9�*�?�';:ZËF�3$����Vܙ��kE�{�N���0u�\k|aT��3G���"��y�S�yH��"J�A��S+HE���2Rip�m~|����� �ܰ�a\Y����+���LQ�l0��F��j#w���	(���B��Zx�.���E� )�&/PP���I̞��>�h�5,Wlr�r%)cA�]���7'�Ћ�l�T�(��ԋT��xB{:i�2"�,�>E����\�vś��Z1`�N�ǁ�f�T���j����k
�ڃB3$�#��]I�r�����n�A8��w7�|��5����`KW����vcy��j
c�!�`�(i3�b9���S�nU�&u������P:�UT�P>&�&i��w��9+���Y����������Z6���E����F}�=Ll�����,۽���dט�w��QP��=2������}&d�X0�� ���3�ҺIÙ=�H�S�yH��"J�A��S+�:G�W]�5����`Kf��}u�귈nIg�R���]6���b9���P9b���dט�w���%=��ބ�����}>p~z�r,J����!_�IÙ=�HB�q;�~ ?�4��ic�n쯎+�ܼ�P����Z�j-J���\�v���GAџVp�m~|�֩������/�-�o%Ǩ��]6��l0��F��j�mV��5f�P4ǲ `6&��Vv�9gP�U,�2������}6S������zL͊�q��應�y�SI��'�����1H}�ɐ��/�W�A�&hH\JHn��z���o�K���g�,P�n��
��D&e�2l��4�y��ɦ�@^7&ģM�'n�^0o�<:�W�_ĵn(���˧�0z�cULjaGkƊ~F˯�+)�"j���b7|#9���hY����r�{p7�j�pܔp�l
d�o�R�GI$��ǂcY�~�s<��MR�������c�A�L'G~��6�7�5�%]���a(􆿳�ټ*w2�56�5����`K��M���o�G�m�?�~ǲ�`�'n�^0o4��t-s�I��RhF��2|9��p�m~|���\��j��<%�a���k�79�����\�vŜ�H�伭�m��3��p���H����Q#�?���;���N�C��{�I��'��R<�����á�~O�
[/��̟vzL͊�q��C.W26K�~�J�� m�������.��R�}vJ^A"�=�f!���)��� � �����p>��u��>п�p=	�˳͠m�xW��9u$d9��}ϔ���GS�����n���㬺ƃ
ᾆ�x�T�\ ��`��K Y�Ћ�l�T�Q��O�بeD�I�1#��Z�����XP���#���1���Q��ǺΕ}a�/�kj�O7��@ׇ5����`KVkLs��dJ�+���LQ��b9���Ȓ��u׿j�h�<��p��޸w�J�W��7/�]�N��&�}c��ko#a��|%G�]�!��	Ǹ�y85���t[�L�a\Y����+���LQ��2���O�}��M�+�'�̗�����C�M�����T�\ ��i3�|)sՀ]�N��&�}c��ko#S0,H�2�]�!��	Ǹ�y85���t[�L�a\Y����+���LQ��2���O�}��M�+�'�̗�����C�M�����T�\ ��i3�|)sՀ]�N��&�[��m�Ua��|%G�]�!��	Ǹ�y85���t[�L�a\Y����+���LQ��2���O�}��M�+�'�̗�����C�M�����T�\ ��i3�|)sՀ]�N��&�[��m�US0,H�2�]�!��	Ǹ�y85���t[�L�a\Y����+���LQ��2���O�}��M�+�'�̗�����C�M�����T�\ ��i3�|)sՀ]�N��&�[��m�UȞm�2GS��a�x�����7���{r��K-��:c_]�8���/����,D�K��D��`�6�\�f��E����F��
��D&e�2l��4��a��se�ξ���I��RhF��?�1�{}�
�?��V5VM�d��P=�<��p8�(�E;*�}Ւ�~ܔp�l
d�R�.��On��M����A�m�(�Jٯ�n
�
�CӞD!�|_@��0�-�`~ ���􇃬Tk��A3�(N��㎏qló��@d��שI4��欱���j���h�߆��y�����DzL�ł)w��������yxZ��j�
����d�R�wX��}�
�?�Tq��A��s��tcb�A���+�J��Y�{'%s��.|Z���׮	��48ܼ�P���MN�-���8���/����,D��8^a�F~+E��XQ�$�E����F��
��D&e�2l��4��a��se�ξ���'�̗������� >��Tb!��u�ϟ��7�4�.1p�Y,�}�CU�+v�rs�i�qt� +�,�T:5�����2������}°������R�wX�ո@����gG���:���U��[��c��w��z䮃�0z�cUL��9v�������ff���-A�¤�x.�Knq���;W��ZLN�	��HfS��1�w�<om����եWT�.JVW{�-v���m��3��p���H������7Pr��ġ��,�~,ǽ��D�P�E6�ټ*w2�56�
�CӞD��VU[��1�
������H>+�w�\w��0]b!��u�)���A7��M������Q]� _ό���.� ��h��UJ�T�G���
�
��(�&��Q�r�rs�i��9˹$m��U2��53��Rx+*H�p�.Cf�����`DPߺL��`y���h}Nw�����k~#���]�!����w�Հ�x9���7�l�|�x �'���XwI����"�]�N��&�G9�:Q���u��N�v{AԢ�a\�D�����R�`�|��K�z�H�MPq6.�T�\ ��i3�|)sՀ]�N��&�G9�:Q��?�1���AԢ�a\�D�����R�`�|��K�z���k��$a(􆿳���2����.JL���Z'h�	�i^䖬n���ȵ�ixUS�D�����R�`�|��K�z�H�MPq6.�T�\ ������q�f@��L���N�b�'Be����s:�L�6yd(7s�9���on�-�6��
�jW��D���M���o�G�m�?�5:�7�+p�R<�����á�~O��L;Л��|#9���b!��u��Ɔ �����Vd�!�`�(i3������� �����p՚��l��Hr�<Uee���R�}vJ^�9���x�����,DTc�~y��i����u_!�`�(i3"�,�>E���]�!��M8���	D%��_�ͅ��r�&U������G|M�#ã�fޅ������ϲ�CyW�f�tR�wX��}�
�?�b8IU_h�΁�a�n��!�`�(i3W���D��g����H���	N^�U{xN��i>r�<Uee���R�}vJ^2nq{�HQ�}�
�?�N��	�Ȓme":l�n!�`�(i3��lJ��튝�b�Bϱ��R<�����á�~O��L;Л��|#9���b!��u��Ɔ ����6���!�`�(i3���+�J��Y�{'%s�h�v��[�x�X���+���LQ���"X��[��Q[R�7ݓ��E�/�����	��c5'!�`�(i3ғ�vq������T�=�;^�6#9���k��$a(􆿳���2����.)}���/��C�x!�H����0pJ\�!�`�(i3�n`5�fK��0z�cUL3�X�j�{q����'6���;8=�g��U-�e���b P]��i�"���$���5N���@^7&ģM�'n�^0o�<:�W�_�l�J;�RQ�y�� Y{q����'6���;8=�g��U-�e,%�0g�����L���N�b�'Beͧ��&�~L!�`�(i3�[�l\���$����b�m��,���b�U�J޿�ġ��,-+��B�Gݓ��E�/�����sc�̆�!Ym��q,�D<�7��V�����T�=�;^�6#9���k��$a(􆿳���2����.)}���/��C�x!�H���J��Ӊ�,�O�%p���ĕ\�AԢ�a\蟖�S� ?�0��E|�,°������Г�����aZ��qA�ETc�~y��i�v1a{J���ǔ���� >��H�݁.�q�-t�A�ݧV��
fJ�	�LÆ���#���x|qj0�ҹ���+F���d���'/�)�ep�d�٣���������ݹ�0���f�Nd+l��p��;z���$Ι��o;�¬pX��g��U-�e,%�0g��հ	�A��ԡ�}s�Z�|�i2C�D�]�!��M8���	D%��_�ͅ���(��ԋT�<����*�כ��p���lC��U�T�\ ��[�ǈ������w`qԴ�~`����vQ� ��}�
�?����PE�K����/�sLgwe�ŉm�m�jp=�>��o�
�v�ξ���C
2��>�o�9�1�Z���=��L;Л��|#9�����\�I�N�_V�ܔp�l
d�o�R�GI$��ǂcY�~�s<��MR�������c�A�L'�O�({������k��$a(􆿳���2����.C�C�~�N���$��R�lDb���(p�+��t��[r]Q�I�������!3ةI4��欱���j���%���3�!�r�A�N!�]fu�Z��"R�bK�s�} Oag����W{~��=����;��krk���:�a��Y�{'%s�[�&B�踫g(�r�2������"�*o�yG�qڒH[91�Z���=��L;Л��|#9����c�hm�i��f��;Z#����n�4�c_����+#��.X���*"v%)��Qcm h�]�!��	Ǹ�y85��p#�j\1�Z���=��L;Л��|#9���b!��u፞�f
t斃���n���g����Qe�2����&���Z02��<��Y����}J�|���|���I��j���S�����0p��t-߱�~����Lu�G{;��Tb����-9�,��Ln+��<�I����,٩G������F�DMs���{��Ń��Hm����AU&���#������`X��{�j�e8�W{4K�)s"���݇�T%{�;����f�kN�ı*�7`����\Z��K���^���?���5����`K�g��&d�X0��!�`�(i3JHn��z��x�f7﹏!�`�(i3!�`�(i3ݻ��A�I4��欱���j�����r%����m��3��p���H����Q#�?���;���N�C��{�I��'�]h�(NAP�~@�\��"�,�>E���}�+�r1D��y��nv�@�ԩH��٪��(2�a+z�K� j��������n7,�
��b3�����>��2��g��@�OW��:I��'�]h�(NAP/i�\	t��Ğ�����}�+�r1D��y��nv�@�ԩH��٪��\N	�����ߦ ��=(!+�C�r�X�pǓ#5����m��3��p���H������7Pr��ġ��,5��=XI��'�Õz����sY?�g>�E����Fy�ӓ��Dc4Ƥ ��`�z��Y��),�B۸�`s- �'|�����:'�>����߰rE%�6��IG��&1����S�ݣ:�T��;�Z-@k�%V"��ߜ�*�l8�b(��+�w]�B׿�ġ��,�]���7'r��VYW\W���}���i�������Z�����9�!�`�(i3!�`�(i3!�`�(i3!�`�(i3������U!��� 9�n�?�����C�G���-��(�O?!A*�7`����\Z��K�����ޣ�bL}b����r��-�W.���^��\i�@^7&ģM�'n�^0o�<:�W�_ĵn(���˧�0z�cUL�_��._0��y	����F��،°������R�wX��KM���d��7Syv�J�Բ�����D�:�d�>п�p=	�˳͠m�xW��9u$d9��}ϔ��F<�'a��Tv�@[�JJ1��P�M���L;Л��|#9�����:�<�L�E��w*e�΢���v��|����OxtX+�Y�z�**ߜ�*�l8�b(��+�w]�B׿�ġ��,���}���7�]�!��	Ǹ�y85�9)e�AjL�E��w*�t%��zxa(􆿳��?ƾ�s��	��6h��LwN��6�o$�VXc_����+�˂߮<u}����Tf���-A�¤�x.�Knq	6�q�i�d�<om���h�p�x�ɧ�	tc�����-�7Syv�Jы�^�)��"X��[��Q[R�7�w�>��p�&���A�&�ʜ���JT؛>�a�W+`�x�oP��@t�&�e�5
���7n�׊�p�&���A����!@ʛ��RY��Ɛ�<["��+�O�G!s��y���S)@^7&ģM�'n�^0o�<:�W�_�܂+�: �mh��LwN��6�o$�VX/��q�&.������Hb�2�ǏTDZ��O$�E����Fv�@[�JJ혮��ר{lGD�V�Bf�Nd+l�Yҽ֗��i�ܰAb!��u�d��}U؄�k]m��¡J���a�GYs��$;��H��,x,����ar�<Uee�N�����H�OM��`�@����gG�x���يj}c��ko#�`F�_2���X�o�!���	����}q?H^��2踫g(�r�N�ǁ�f�TpD��ZOU�ό�]2.������Hb�2�Ǐ��Pn<����U�9*�v�@[�JJ�-t�A�݆�ŋ�R����@d��שI4��欱���j���-+��B�G}ϼ 8���hy�`�w��v1a{J��~z��k�Ɛ�<["��+�O�G!s��{lGD�V�Bf�Nd+l�Yҽ֗��i�ܰAb!��u��@��A���k]m��!�`�(i3GYs��$;��H��,x,����ar�<Uee�N�����H�OM��`�@����gG�x���يj[��m�U�D�d��k��X�o�!���	����}q?H^��2踫g(�r�N�ǁ�f�TpD��ZOUi3�|)sՀ��{�j��+�g�>U�wE���Ov@)�l��0�L�E��w*$��O�&���f�kN�ı*�7`����\Z��K���^���?��5�e`��9����V�,�Z-�=�"�,�>E��Ɛ�<["��+�O�G!s���bl�_�p�ξ���I��RhF���k��76����,D�ʥ��G�Q|�P��Ȓ�0^M�U�î�D�p�&���A�&�ʜ��M�l8�	
ڶ�@d��שI4��欱���j���-+��B�G5�e`��9����V���V�%�1��9�29jƐ�<["���܁�_�jZ"]�Vp踫g(�r�N�ǁ�f�TpD��ZOUi3�|)sՀ�)׺������Y�U��3Y��P4������jL�E��w*e�p�������
��M����A�m�([}�@��L}�
�?��V��G F��x�������b�W�[r��-�W.��@��i�=�f�kN�ı*�7`����\Z��K��4����/�Ӝ�z@����U��@at3Y��P4������	�v�@[�JJ혮��ר�bl�_�p�ξ���I��RhF���k��76����,D�ʥ��G����9�~���&�����Q]� _�� ����/?(��=՜r�<Uee�N�����H�OM��`�@����gG"�t�'ێ��0+��?�z0�塴`�n`5�fK�gh1�͖5�Zz2|��M����A�m�([}�@��L}�
�?��V��G !]�~F��A��yU� �7s�9���o×��̙�F�9 }�m�f�Nd+l�Yҽ֗��i�ܰAb!��u�zk�����>�P,љII	��G)��d�٣����Qq�M��H�_�ЩI4��欱���j���-+��B�G�����bpA���3A�Q���jμ�Og:Ba=�d�٣����Qq�M��H�_�ЩI4��欱���j���-+��B�G�����bpA���3A�Q���jμ�FJ���-w��z䮃gh1�͖5�Zz2|��M����A�m�([}�@��L}�
�?�af��pD�Ї�6~���^���-��b�W�[r��-�W.��@��i�=�f�kN�ı*�7`����\Z��K��4����/��)}���/����ly�P�r��n�Ŀh.�wK��� v�@[�JJ혮��ר�bl�_�p�ξ���I��RhF���k��76����,Dv�	}x'��֢��s�K�^���-��U�î�D�p�&���A��J2N��{lGD�V�Bf�Nd+l�Yҽ֗��i�ܰAb!��u�t�,�NL}�="��x8I���]�q�GYs��$;��H��,���E���:��`�z��Y��),�B۸��L� s�j8Q&ֳ��eew���m��@oX�� Y�]�7Syv�J�Բ������sl����?r�<Uee�N�����H�OM��`�@����gGdR��Ƈ�r��F�f�J�㴭+�J��X�o�!���	����}M�l8�	
ڶ�@d��שI4��欱���j���)@����Sb!��u�d��}U؄�k]m����!怬��L�E��w*e�p�������
��M����A�m�([}�@��L}�
�?�^)�G�B�+�WdM4@��CX�y7Syv�J�Բ������sl����?r�<Uee�N�����H�OM��`�@����gG�x���يj}c��ko#�v�W�0�v�@[�JJ혮��ר�bl�_�p�ξ���I��RhF���k��76����,D�x�/��Y#ѥh����܎�Ɛ�<["���܁�_�jZ"]�Vp踫g(�r�N�ǁ�f�TpD��ZOU����q�f@rD�9���S⏸[����Q]� _�rs�i��@�N3,(�;^�6#9���k��$a(􆿳���2����.�N��+�j����tL�\�7.��Z鎬�������(����S� ?�0��E|�,°������R�wX��}�
�?����Н������\d�7s�9���o��S8����ٺ?�n���㬺ƃ
ᾆ�x�T�\ ��i3�|)sՀa�K��U�_3GH�F���YD���xZ鎬�������(����S� ?�0��E|�,°������R�wX��N>�4�
��o�M���]���!E�.tik&�#�Bp��!�ʆ�In��tw�?�b�>޼�\�v�	�+�&I(&�L����6�{�Pe�E"���m�PU��i�2���#M*�1̞��>�/=T��?�N���������!�����T%wxE���8�V����8��?�d���&��뷖iU��5i^��pn��^��(���B���Q��ǺΕR'),��`��͐�4�E5$f��_Ub���uQL+��槑��gL��dn��A3��0����$��Xo����Ǳg�P�e�9؏�	���ul0��F��j�.�p�2�z�����������z�'Ty	��)~�W����1�S��*�7`����\Z��K�����e=_����開�E��ч¼xE���8�|`��P��2�;��	1�jݭ�F���E���%�a�<�W�C%��p��:յ[+8��x���	R����>�ROQ�U�"��>��x2���y]/�qF���V]��y���KT��$E��	��x������a�"�i�_:���
��vK����0/ܤ�(g��V�-4�{>���5ߧE4��?�{�XԪ��]^)��������w�s��q!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3���aR��$��Xo����ǕGF��a�1�Z���=�Ln��S�W�.�p�2�z�����޴�ik]�_�8V��FU"�
hYY��B�D�F �(����C�EPj�x�Z鎬�������(������t�\~ �g8Yw���k��$a(􆿳�ټ*w2�56�5����`KIR*�fN��/��+l0��F��j�bOM�P�C���_�\G��4�	B45�EOs\�̞��>�nQ�rV",�Ű��dט�w��5kj�Hn��O�z���@��]�h��)w�<�_N��W���-�JP���It�Ɍ+8�3��$<�Q�R�j�`��2�.�05k
��F�2�q#O��*V<�ɔ�,���T�K�TZLk]�V�Y�\Jm�A���(���d0J�̛�ĭms)������*��?���-)zd70ǰ�5aj�r�[�"�@��e���ú��'��X�T��A���sG�]b�` ���"�+�*�p�a=}���dm���lD��~��~�
�b!��u��D����e���b���Q]� _�rs�i��d�	�6%�����ׄ����ӯIJ ��`y����@����gGD=�^�(|���Y�ǒзq8�Ј'���Xw���,D�Z5��جl�l"���E����FZ鎬�����
!-�n[�=�5x�=�C��Y��]�!��	Ǹ�y85�����څ��;�¬pX��g��U-�e,%�0g���[�=�5x��-�f��_�]�!��	Ǹ�y85��L�@��f����k��$A�h��+Fen����9��0|~�LL�a(􆿳�ټ*w2�56ݓ��E�����aGl���lJ��튝�b�Bϱ���w�K�1c+����Y~�y����u{ᵿ�����"X��[��Q[R�7ݓ��E�S���%���lUR^�p��b�Bϱ���w�K�1c+����Y~�y����u{ᵿ�����"X��[��Q[R�7�׎o�|䖬n�����lJ��튝�b�Bϱ���w�K�̄�Bq���ZLN�	�����#oM|#9���b!��u��d�@���GL�q��j<�AԢ�a\��F�dH��|c_�m��ġ��,�z���a�R�wX��}�
�?������3�� n��P"G�wk�١��	;q}u6��\����m��3��p���H���F`���G���`y����@����gG�' ��&-,j%b�HۭxZ��j�
�iB{�Z�_���}�\���0�=<MW�-}�	mp�?IK��y�8���/����,DJΌ�#<����Gq��T�ٮ|�,
���1��e0����yN��7��aq���E���ss�T�\ ��i3�|)sՀ/��{��`��NۥUn�cq�����f���,(���B�����(�犽{Tɀ��k�V\���"X��[�w�����@����gG�0����O������Z鎬������_�,�;�7���c��չ�Ad��d�٣���N N�S�qg2�K?\�E��ȷ���n`5�fK�\w��0]b!��u�z�
1���;���+�J��Y�{'%s��jb��:0�g��cH�wA�?�*42�����`y���h}Nw������S�зq8�Ј'���Xw���,DU�m#j[����L ����b�Bϱ��ᵉ3���P<t8��3����開�{�&�;G�<t��Et�{Mq��JG�4W��(�!�>��y�P}��O��ꅽ52�����8-|�D<���K<�%�/��Z>L�<��˓��>�X6�j~H�RtV�^������h�g��cH�wA�?ܣ#�'a�������2������}�ޥ�6���Cn��P)�A`�>;�;F+W���F�^��NPSI�-6��f���-A�¤�x.�Knq��H�����ġ��,d��^��H����8��?/�1�8fÁ��/�6�£wO��l��b}*�ZLN�	��!��"� +}���k$ �����a�"g�]@n_���?3�j�O����9j.�l>'�o��&LI |���\bU2��53���6��������_�\G�k�y'��aum��x��m��3��p���H����HRCJ��<om��'@�(��P�?�R��niR$�Si"HN��R���ء�I�Ǧ�;38K��1X�7�o���N��i�m�ڨ�hծ�5����`K���ػ�T�p~z�r,Ln��S�W�.�p�2�z�C���B��	��u8-�_���Cg#�@����gG�XpAS"Y�j�`M!�`�(i3"�,�>E��P"G�wk�١��	;q�� ��-�BM�ܤm|�8ɂ�T�T�\ ��i3�|)sՀ;�7���c�����-ќv���z�Ji�!�`�(i3q��T�ٮ|�,
���Z�˙}���.ᬵy��"C�����T�\ ��i3�|)sՀ�`&�;y!�<����i"��!�`�(i3±�sR�{F�{xy�b!��u�v�A�
^^3�V�C��k�HvL)���(���G
'���Xw���,D�8���Q׆��p0�Ĝ(�IyI �q�T�*�u��6�\w��0]b!��u�v�A�
^^3�V�C��k�HvL)���M[�S���]�!����w�Հ�JX-�ܶ�0l�x����b�'Be�s�r��<��n`5�fK��0z�cULA6{'8�0��9gP�U,�2������}°������R�wX��}�
�?�&aD�4�X�X�>c�.A�/v�K7%'�d�٣��c�A�L'����8?�o[L��h �=�.�v�L#�?��Q[R�7�n~�x��Nh���W<˥�'ܤ",Ц�} m�g�z�&��Z鎬�������(���_G3w�
|:
@�!]�������d�g��U-�e,%�0g���JX-�ܶ�0l�x���
��e��a�����!�`�(i3�d�٣����Qq�M��H�_�ЩI4��欱���j���-+��B�G�n~�x��Nh���W<˥�'ܤ",�X�G[�/v�K7%'���+�J��Y�{'%s���gt�͓�ξ���I��RhF���k��76����,D�8���Q׆��p0~�5�H��s��ꮂ!�`�(i3�d�٣����Qq�M��H�_�ЩI4��欱���j���-+��B�G�@����gG���U�\ʭB��2�k1�h�H��*F7	G�<�*�P�ߚ�6�xZ��j�
�iB{�Z�_���}�\���0�=<MW�-}�	mp,��_А#�<om��]T����?�T�\ ��i3�|)sՀ�)׺����\� C&����q��Z��2Q�g)/�_~�:N��n`5�fK�\w��0]b!��u�q���3��`��R�`��ƍ ��_~�:N��E����FZ鎬�������(����`(�WOݥ��{)�h �=���"X��[��Q[R�75�e`��9����dz����NR�p�'q�-��nEg�N>Zh~dTfX���b�Bϱ���w�K���1`��vߜ�*�l8�b(������l__�I����J�����g���R�wX��}�
�?�u����p�����+X��FJ���-�� �]q"�,�>E���]�!����w�Հ�b02�O�0�5G,��Gc#%@Ԫ�!�`�(i3��Q]� _�rs�i�M�����geE�vx���ƚP�& 5f��e�T�\ ��i3�|)sՀ��K���B�V�C��k����?dq���z����7��,��S��]�!����w�Հ�j�|�{'�X�X�>M�a���;}`O�k�
�p�	%6�d�٣��c�A�L'��$;-,�J�d�@q�2������}°������R�wX�Ֆz�6�g�u�(��l�/�沣�*G^+�(���G�����}��e�C�q�뢗�˯��Wނo̒.�9�lA���k3����)׺����\� C&����q��Z��V�X8�9a/v�K7%'�n`5�fK�gh1�͖5�Zz2|��M����A�m�([}�@��L}�
�?�u����p�����+X��FJ���-Yk��P(I"�,�>E���]�!��[@�zZ��g�f�kN�ı*�7`����\Z��K��4����/���>��왩�/Tu����W`GU�!i&G�\��u���9�9�ƭLF����� ����/?(��=՜r�<Uee�N�����H�OM��`�ȓ�iӚ/2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hCݮ2����g?mЛR>2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!�V��2�ќh~-s/�{pў�%63:��ۜ���=0���m?�>��?�%<h*\�J)0�	J���j/ǈb��
J���%~k�b��W�FzFp�]�j�
,Z͚��Wᜈ��� C�_�Z��`D�EcX1)!w�G37)ǝ�,^aj�+��+-2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�����z�}�+5�4��c�.}�uP����}�t콢��0��d�@����i7N�_�z*K��I4��欱���j����Eo(d�J��:�����`�x���I�?g�f��Qө}�8o�C���7I���ʚt�  ",�PM�^-q�x�l��1:�N�*�xS�_�p��á�~O���-@t�/�W/S��8(�E���Kt�K��^��b̞��>�h�5,Wlr�r%)cA�a��OY��]V�H7'�R�^Ƒ���)ύ^��R�^Ƒ��f�?ǉ�=�]{��_G�D�� ��ۋ�/�ͪ!�`�(i3C��[�����p��@LC��[����r%Ĵh����ڃ�"��
!�7��}���3r�e����kn4@Q�/�!�`�(i3̲�2�!�vc]x� ��2[QvA���^à�١w��zj~�X����>6�b N��t��f�?ǉ�=�[b�0<�Ԣ�{��W�����A@�
�s�?V��j�c��<n�p�ϟ��7�4X�֐�._�ݚ�Н�l��A-���:��]]t|��sQ�G���+����rV���qޤos�em������`��B�'��a�F�,�U6�Q�L��
�:qEp �D�lh8t����sV��o5]��hЗ
H�ǅ��$���F���:3�U�;���N�q��Xr�;��|B���r����T 3���䟳��L��C����N�ǁ�f�TpD��ZOU_��s�֙7�}�!��P� d�c�m�/N0
���U��G)+��T�����D3���t�  ",��ݚ�Н�R�7h�,b0V�u�Q�ݚ�Н�¥������]n��-��w¹��<d�,��L��!�`�(i3��.��֞�������i��D��;jQ�#���F�;�@"��ݚ�Н����8��T�h���}둮j\����C��rR#K�p�ݚ�Н��K�^��Q��G�S>\.�!::tm�0�i.�9!�`�(i3�2*Q=F���q/���<�����7
!�`�(i3�dv��oTN֢&@��&!�`�(i3k/�z�xEQ���*[UxG!�`�(i3��|��p��PIQ#�C,0�?���!�`�(i3��9��稕�a�/!O�f�?ǉ�=�2��}��CϾH�)�V5VM�d��m�.j	f�?ǉ�=�2��}���zgm##��V5VM�d6��0]�1�v�9�ʅ.�g3Z�Ǵݵ���pÓ�}<�ž_�F�Tq��A��s&?Z�l�(�u��@t�qP�V>tI��RhF����u�*��?�d���&��ݚ�Н��V5VM�d6��0]�1�g�)�I��#�r��8��ҥ�|HN��R��?�d���&�Tq��A��s&?Z�l�(�����0`;�V&S�b6j�"Hsކl9�p������l��Vj�Ra�m�,�*��'��ҙ����
�Z�S$J�	�LÆ�c�9ʼ��$l'>����J��:����9�{�Jj3�a�5@�i�QR�j4gM�+5�4��c�� D�_\HN��R��?�d���&�+r�^4Y�BM�e�x�U3u��� ;��|B�.y7bژIl���o���8�:�����zV���z%�/��Z>L�'��D(M&��w>��Y��$1&O� �k�3��6J�Ko��ih�|����
�Z�S$J�	�LÆ�c�9ʼ��$m#�P�J��:����P� d�c�.1p�Y,��J��ۍb�o��_�Rv�䩲$����tb�����+�^n=\f�5>����Db^�.1p�Y,0Y�X��f�\���F�`yx�>�+X�M?��y�!�`�(i3P���x�NS���U��[��c��3|v��Eb�z'hۉ)��d�7�q�՝� s�#0�ʂ�j�Ï��	�l�lM�3 H�RtV�^�s�Yls��8��GM��-����!�`�(i3P���x�NS���U��[��c��5H)�c�8Qł)w������U+��_����E�ł)w������U+��_ �2��9gUS����a$�/ϟ��7�4�.1p�Y,+
���Q�"���Urܰ#y���:5A��pfĉ>99��A0ok��fĉ>99��A0ok��W?�;�끓��~�Ly�$�|�m��Z�f�WM8}�	76�&�;��|B�mC�8	�XB�����C�����tP��b&�\JG8q.j<��IZ��x�,y�#���F�F��b�\��Se���7�}�!���V5VM�dC��6�g����5�ź�+���*#nC��6�g����5�źP�?v�l��+�ϸ�i���U_&�W\�a|��sQ�G�3��ݹ�w5���i�w�R���y>��yСQ=!�e���26}�i���:I�#��y�$�|�m��=�_�7V�o��_�Rv�䩲$��GQЌJ
��`���φ��<�6��ߙ�[�>	ol�~{�Ž\���F�`yx�>�+X�M?��y�!�`�(i3��6J�Ko�����P��nF���<�W�.�P�	��
�Q�}�k��^�1��dc�@c�����h��-����;�jmT�#�,l����M?��y�!�`�(i3�<��7gҠ�(�2ʛ[�q�ܦ	&�P��k�Ӿ]ܦ	&�P��UB�I'9gUS����a$�/ϟ��7�4�.1p�Y,v�)�DZ�ϟ��7�4�.1p�Y,Q� R��F}v���۹�
�:qEp�;�P�t�5fĉ>99��A0ok�׹�����A�;�����[�F$�kj���6J�Ko���zX��-Z�+�ϸ�i$x���z*�7`����\Z��K��rt=ٝ��b&�\JG8�j(&
M�K�<�
�d�ξ���'�̗����
�t�c��5�O�%E#Pc�{��lq�<b*�_���t�T��?E-h��`f���s��6}���iI9�o«IX0F�M��6J�Ko��hm�ko@h�H����Qw�c4~Nr_�mS8<�n�ݚ�Н���� ff��X	n�ɺb_X�XV�b�z'hۉ)��d�7�q�՝� s�#0�ʂ�j�Ï��	�l�lM�3 H�RtV�^�s�Yls��8��GM�`�(�4�bł)w������U+��_����E�ł)w������U+��_ �2�Ъ��tj/�՚�-����!�`�(i3�<��7Nǌq�p�IC&��b��mf-W�c��ǳ��&�!�`�(i3�5ߧE4��!�`�(i3�5ߧE4�퉅�%>�rG߸��S�Ȍ� �Q$j�sP��':�HN��R��?�d���&�x�����<����՜����� ff��pH�x��]'\gWg��	�Z�kfc?�#	*]]�iI9�o«IX0F�MG�k�P[�;�jmT�#bs��2[�a��o���H�RtV�^P���x�NSB���j%Ř�I4��欱���j��������my$�N��o�/���;�Ra])n#���^a�nu4Bޗ��jw�	���ݚ�Н�y�}�6f&r#o�]�ʄ�lZ#s��kgҠ�(�2j�y�`CrgҠ�(�2L���yF��G��Hb� h�ҩ�,��G��z#�r��8ߞQ���l�N�����K����F?Tq��A��ske��|ξ?�R��n�#ٷ�Ef��ݚ�Н����F��O��;b�-�2��;�P�t�5W?�;���z��O�Q��D��y�t����M~V��	��y��E��D�VvA#&��Q��r��`�@2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�_L�oe��Em�Ԣ�+d%�4.P�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcN�H"����H��X�����k楊HaU$kX�M�ŗ\�'	�?��[n8�A�A���p������'HY-��Yk"1/|sL'���oֲ󄰊�t�  ",�PM�^-q�x�l��1:�N�*�x�i�ۑ ��GZ>.�0�<P��C���U��+�Xa�H(�˕,���9^-��w,�����<v���G�kޮ��n���㬺j;��q,9��n�7�Y����X1Ο<������.��R�}vJ^Z_V�`��n�����������_-�ȩ:T�v��1���5Z��L/���?T�x~1�@����Ի��= ��j���}9s�X���@�X�ƭ�i�\�;�WQ�.p�2������}�k�+9=��X�u��
)\Y����i�\�f�~�ڳkԜ93�����U�6n�jD�pϓpy%����ڻ�<i���eŞuT ��>��p����nZ���t��˳3[�u8��⒍~���*IϢ���z>�6����iA'R�	�2�O
�� �ݚ�Н�+��%�k<r�`�ab8IU_h�7��m�K��ݚ�Н�0q���Q�L���/��@��e:$h�7�cl.�	�C�
�:qEp3?���*�k-r;�g�~��nސ��W�`=#�eH���%�#�o����q,� L���门:<#�'	�?��[7�}�!���_fy�:�K���~�����G�٘����������)2��V|j=�����.�8�������0�Vn}�R*�V�K^c�{����]�'�g.J/-�����H��2�6.FwZNEߚ�/{j���혅vº��H�:��a=��Y��),�B۸��8�B���ow_;O
�J��:����-��ټsU6гdP!3)T�ϟ��7�4K�ǟ
��)�;b�-�2�V��	��yv�ʯʗ��/{j�䰜�}Dq�f���t���R��4�|W-���Y��)�D�YG�9E�g�������(ӈ���m�r�����nސ�ш�A_�u�x�y�Zgl-�g�"�����yb�z'hۉ)��d�7�qą.�g3Z�)V��B�1*�-�!�/��P�	�#ʁ��
O�߰�b��v{7!I���6�{�Pe�E"��*X��[��7%^�W+��W�}�
�?�G��-�HG($R�i�Yl-�y9C�M�Y�{'%s�h�v���j(2z�ܼ�P���MN�-���8���/���}Dq�f��
�CӞD��m�q�/�Wv�A���n`5�fK�\w��0]"(<K�'P�1r���!�P�)��xuo��*h�/^!���Z鎬�������(���b�	�/ω�HM���#ga(􆿳�����r9E������y�(����<mG��-�HG($R�i�Yl-��8.���B�Ы0�Y�C�x!�H�'�İ!��eA{��'�K����k$ !�`�(i3!�`�(i3��7I��ٜ�}Dq�f���ŊPT��b��Bg<���P�5]'\gWg��	�Z�kfc&�2����{y����i�q,?5q��7���9�:)�
�9P/�%��F��H����Qw�c4~Nr_�mS8<�n�ݚ�Н��T�T�y�8�Hj\��9��T�&�{_8�Y��=�}�Vݨ��}Dq�f�c�{��lq�!�P�)��xuo��*a���P7��{_8�Y��=�}�Vݨ��}Dq�f��k��^�1��dc�@c�����h��-����!�`�(i3L�J)���� \L�1tSjv�!�`�(i3G��-�HG($R�i�Yl-���^���m�q�/���e���W����^dE���b��Bg����;?9gUS����a$�/��j�4�<�..�4�ᜯ}Dq�f�Dw\���B���Q���X��+M�j�/l��I�mۯ��uz���O9�(UҔ����F릴�˼�RZ��P�k��!B>gX��کb�b�������Cҷ��e�A*�����b��Bg|:�X]�Y{�<�������̿}v���۹�!�`�(i3���F��O��ݚ�Н����F��O��;b�-�2�$�)�vx���Db^�Y{�<����
�9�vm�ڨ�hծ����ҧ� 4� I�;��wñ�_
���.{Π��yGb�:"�G�}��$1&O!�`�(i3�Ե����d�φ��jp�m~|�֢�����k5�D7�B�'��a���L�jA��h�5,Wl�/�O'�=��8�Pz��Z鎬�������(���/%Z�ڄ^1JK�2$�h"x�����F��%�>&�&i��B��9�OG��-�HG($R�i�Yl-%�z(�~�:)�
�9��3�����1{&��� �A
i�eL!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�{_8�Y��=�}�Vݨ��}Dq�f�w��'�L�����P-�k�+�ϸ�i
9'�@@��!�`�(i3�ݚ�Н�<�V�QK�}ܱ������١@��R'cf���³5��*�7`����\Z��K��qb	��G��W+��W�L��@�a��<	: �v ���\{H���7Әi��7u�`��Y��),�B۸�Үo7�hm�ڨ�hծ���%>�rG6j�"Hs�07�)(�~��k�u&����A@ž_�F�w�R���y_Nr`e���f��*��]�]V�M�ujVA�ڦ�c42m�O��{��;Ӝ�+:�h��"];�.�� �\�O0U'?�d���&��ݚ�Н�b8IU_h�U���H^���R�}vJ^&�)~~;dN�<@Iv��nt=:��:5A��pt�td���5FwZNE�����A@�����	�+5�4��c���s��1�y�n�F�:)�
�9f�!�Wm���m�q�/���e���Wƈ��hZ?�JF!��D�����k$ !�`�(i3!�`�(i3.�`��ai�t�3���B���KOK�I��RhF��?�1�{�ݚ�Н��,��	r�-�y�4*$�*�7`����\Z��K��	�v�Uū��?�ؖt/�u��]��8�; �ì��O9�(UҔ����F릴�˼�RZ��P�k��!B>gX��کb��l���-0i.1�C�my$�N��o�/���;V�Ո��!�|_@��0Ï�6]S*��C�M$�ѦY�Nj�{_8�Y��=�}�Vݨ��}Dq�f�)�{6�U��'�U$��Y��'���S�[�����E��'Z*)������oF~�S?�d���&��ݚ�Н�w�.Y�[�O��h�|2;$�J�$�* a��C�M$���vdRɅ�tCsd�h���Z��!�`�(i3FwZNE�����A@�>�暩�͚+5�4��c�� D�_\!�`�(i3�.�g3Z�j5�{�=���� ��,Cb���fĉ>99��;��|B������{�X�&����4C"1v�ݚ�Н�<�V�QK�}ܱ������١@��R'cf���³5��*�7`����\Z��K��oaF��!�W+��W�L��@�a��<	: �v ���\{H���7Әi��7u�`��Y��),�B۸�Үo7�hm�ڨ�hծ���%>�rG6j�"Hs�07�)(�~��k�u&����A@ž_�F�w�R���y_Nr`e���f��*��]�
,O?2@@I��)���W�w��fD�,��ϬL�0v�6���N-Y&yo�qX� �Ĭ1���$L�9���3v��u� 
~�F�,���XF:����k!�M�Z���	�^�̷ؠJ��:����շ���������j�Txk^����2��'B{q����'6���;8=D�P�E6�k��q��־�W+��W��G�dE�h�k]m��,�۞��	�����p�?������D�v1a{J���V!��N��:5A��pw�R���ykb>���p�������nSf��շ���⪞mf��EYzȧ���2��'B>&�&i�+#c����nS�3�ǻ��d���!i�B�'��a���L�jA��\�����b8IU_h�'=��!�̫z�����	HN��R��?�d���&��|��Li�8j�H�pHN��R��?�d���&�zY]�埅��!�ٞ�AW9	 6j�"Hs�9'{Z5xls�]�Ĕ��7n)�26���k楊HaU$kX�.SS�Zs�c<�^<�H�W+��W���	�|Jgq�M�4�9�0��L�w�R���y+1����!���Dte��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���������G�٘裣
j ��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 �a ��^�.�)����x���	R����>�R���mK�g+�Vr���J��:������G�٘�#|�4H�(z�1�:�Ω��]	h8��`��(	�t��4ԲcZ7��n	l��Q;�im��ȍry��	^�R@Κ�2���eip���,���C�M$��k�+9=�}9s�X���@�X��״��/^l�Cn��P)�W��7E��nW���`moF˯�+)ƙ���ល��������6%�a�iyV�[R�^Ƒ�ӭ�i�\�>&�&i��&�C�/�����/�U��֜��3uwТ�
�+���LQ�f�?ǉ�=7�;�r��0I� X�1��F�7��YȨQ�?�Q,\ͨ܉p����O,8�ݚ�Н�Gظ0����!�`�(i3t�%�Z?��<�ry^�Y��
�iC!�`�(i3Tl�������l6��\�LtF�!�`�(i3��c�����:��IK��<EOJ�uxm�3���w�@V�@0�u�����d���e�i��H���ݚ�Н��u��g��L�����S�Zq�%�V���٧��z�?�+�p!�wӨj]h�jsrCm�kz�6/M��:;��krk��~Oc՝��t��e7
 G��sg���y[J3�j\{ف(�7���<��Y�(��/�h��L���2?�d���&�x��7��M!+O��]k��o������"O����@��
�����D�Ϩg��U-�e a⣃_B7�}�!���G�6\��foti�J"�nFW�JyS��v�<�$,�۞��	�>�A0_�|�;b�-�2�V��	��y�� �P�qN��v�<�$ߋ����-V��	��yG��Γf���b$�\�U�2����/z*q+6j�"Hs0vZ��ҹ�[�Ʃى�6����O������"��[�Ʃى��+�@t�L�FZ�1ǝ?nQO��B��N�����?�d���&�����7i��p��(�+��T��/o��إ�8p	�rh5���Z=%�ņ`���"�R�7h�,b0V�u�Q�ݚ�Н���M����3��~ �X;p`�f�Nd+lJ�VeSZ3&!�`�(i3Pt�d��R	}�������O9��Q��Q��O�بeD�I��k�+9=:(�I~�����h�Q7!�`�(i3*bL�(Rp~z�r,,���9^-���2��̪U��֜��3�&8�,��w�Iſ�Κes��O!�`�(i3Vx�%L��]n���@�����T�v��1���5Z���ck�7!1�Z���=������uwТ�
�+���LQ�f�?ǉ�=NM(�n��1�Z���=��m�B��dVkLs��dJ�+���LQ�f�?ǉ�=�A�����y������i�-�����m l�o�1#V���<�dv��oTN֢&@��&��|��p�S�o@�����	�;�ݚ�Н�h�'f R�苇��Fe#OOJd֯��
�	?�<�&8�,�g�Hn7�(��wӨj]h��_--���g�_�C�6%���lи{K��n٬|��VC\�2x���ЈH����@�/�MC7z���mp"�o�%�Ucf�9rVu,� �{k�h�+|�c�$�t��R����s+��6�.��6���N-Y&yo�qX� �Ĭ1�z����ْ��4F�;��%YM�	�v�3�2������"�*o�yG�f>x�:	�W+��W�1h#����5��������o��D[�h��4o�ݪ��H��q�/���˚����Z��!�`�(i3��f
t斃�B�ӗ�zjJrf����G�m���*J�X�$����q(	�fI��)���W�w��fDv���k��/9ݦ��.�g3ZE��g�Hb�t]�<Lz�B)/D��Aɶ�;Z�6j�"Hs0vZ��ҹW�`=#�e��}�Q�� �F?P�.!wG��sg嘙�^u�� 
~�F�,���XF:������X`��w{���Z���F%�X����)mSj�Txk^��]��3R��������Vo[���˚����Z��8��;Yv^���d����`"*(�D�pq3�O�̑N�$hF ���M7M�w�ToHA �I��)���W�w��fD��0[��Z���zh�QS��:Z�����nd肈��d3���2��'B>&�&i�+#c����nS�3�ǻ��d���!i-��ټs�}s�Z�|�Z�+Ěʮ����?�b8IU_h�¦�naä��E�i�m}66j�"Hs�ĖYS⪞mf��aT��3G?�d���&�zY]�埅�A���V�d��)�(Qe2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WOtl�܎���~�k��`���7�9 �e�I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�F�I�_
S�.�)����x���	R����>�R���mK�g+�Vr���J��:�����B�����혅vº�w�⽒���M����A�m�(�#W�U��ظ�d���!iR����
w���������q�©�����<�������~s���^��ņ`���"���n	l��Q;�im��ȍry��	S�_�p��á�~O��� g$["! ���t�=�v��*"3���'�C}�A�f��!�`�(i3w¹��<d�Ji�];���W����vcyj;��q,!�`�(i3n�NQa"_�?���C[u��oŹQ!�`�(i3EfVNN{s�ܱ?'�EfVNNaJ �!,��z�_�Б�����Y�M���˻��0y��<�ݚ�Н��dv��oTN֢&@��&`
 ֢��'B�ɏ��]�!��	Ǹ�y85���J�%��}c��ko#ƌ0Q_,�F�dH����y�����/��b��7<Rnnx��m��M��ٌ�RnQ���_A}c��ko#��'�Ѱ���w�K�R he��as�C�G���-�p'�"�hPW���[fS����6s!�`�(i3K�\7}�W,g�%Y��̗0z�cUL�����Y���3���α� �m�Ejۧ���Ɖ`���|�F����A�+�~@�\����F��aQ��T�\ �͚Go���{���3���΂�l/�Q/�F(�@vW4��`�|���eC�����jA��L��)��$3˓8���/�f�?ǉ�=q�\E��0�����~���H)j�]b��Ҧ���!�`�(i3�� ߌ��t��Ҹ<��n<���AV2�Q��ǺΕ�A�m�(mk�6F���f�?ǉ�=4%6� �7D���K^�)��VU[��ͮ�@N���!�`�(i3h�'f R>N0Θ��ݚ�Н��\�LtF��c����ҧ��j� �w�R���y����C��a,5���(�JZ�Vk�;��|B�xX�N�C���P�	�#ʩ�Αo��p2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�-I	�\�'���2�V�e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcu0�I
�K��[�Ʃى��+�@t�L�FZ�1ǝ?nQO��Bm�w���i���Z��@?d�s�8K�I�����S�����:�a��Y�{'%s�[�&B����!3ةI4��欱���j����G�"�-�d�uY�ة�;mQ��8���/��8&���I�f|��Jp0�m����!(��'HY-��Yk"1/]���!E���VG%�4ك��	ቢ��S���� "5�]9��n�7�Y�9ηd��K�=5h+�-��L6C\TF��I��RhF����y�;vN�ݚ�Н�w¹��<d���<
DN�!�`�(i3*bL�(R��u��n��ݚ�Н��z~~�Y_" �g8YwU��֜��3����d]���GF��a�1�Z���=�,���9^-�x�	�2��g�P�e�9���6�Q��xj����R���it	�T!b%�ZV�p����nZ���t��˳3[�u8�̇i�d�?�!�`�(i34�0 L?�p���@Z�_F�k-�!�`�(i3�苇��Fe#OOJd֯��
�	?�<!�`�(i3��&I���m�
��,!q�\E��0�����?~K�Qf���?�ؖt�2�O
�� �ݚ�Н�$���]׽�!�`�(i3
=�2����޴�ik]�\Nͥ���zX� �Ĭ1�<^��0�u"��D5�|أͽgF"?�����	N�ǁ�f�T���j��`����OD5�O�%E#P�F%�X��:*�Ev��&~����w]��m�'6���;8=D�P�E6�k��q��־�W+��W�OV�<��V�nX�p��"_.��45��h��[�~�N���|th1�$�g�;b�-�2�V��	��y�� �P�qN2�W1S�]I��)���W�w��fDbYގEV�+pMhƽ'w�R���y"O���%�\�V��#�$��`eom�.P��K`�J¹��ŲVz��s�q@C�x�>���� �4&Ƒ:2�c<�^<�H�W+��W�3qQ�"���M���R'),��`ތ@�'��|0;��|B���r����}ϼ 8�����?�ؖt�-1Z�����0]AZ鎬����
C��8q��f�kN�ı���}J�|���|���{uJL����Y�7#�xI��;mQ��8���/�ݾ�9J�c(&�L�#%i��{a���~�(����5���&<˴m���q~�i��{voPYӖ�����%kR��������֢&@��&�=�<�1���A��|`��"�X;p`�����Dɵ�p�AJ�e�$J��a�U"��zg��p��I7��-5�B�wj$g-��VkLs��dJ�+���LQ�f�?ǉ�=8��ؤƼm��P���ݪ��	QY��K*�+W���F�^�Y�7#�xI���E��!�`�(i3���0/ܤ�(g��Vt����$�����p�><{ �=�%���$Ȧ�f�!�`�(i3���ȍry��	֭�h��Oo��0��7�X;p`�l.�	�C�!�`�(i3h�'f R!�`�(i3>N0Θ��ݚ�Н��\�LtF�!�`�(i3��c�����:��IK��<?V��j�c>ݣK�6<oC7z����t�f�2E����u_R�^�s}�d!�`�(i3�� ߌ��!�`�(i3^8�]3t��xE���8��j�gg�y���!=.�
a�~~��}H_��i�;��%YM�	�v�3�2������"�*o�yG�f>x�:	�W+��W��F%�X��:*�Ev��&~����wd��~TV�.1�Z���=��#t:0���nS�3�ǻ��d���!i!�`�(i3H���7Ә,�۞��	�K}�*��6|��ŌM�ߌ�LM�a$���|f��I�{�P��HN��R��?�d���&�ۆٗ��NJ�F�}қ~ą.�g3ZE��g�Hb�t]�<Lz��al���t�td���5����,�ǰ�QCT�"�ԩ�V��R{�#_�E��'Z*)�6/��������рӚx�mWᅫw�5�O�%E#PFkH���޴�ik]���7�i�s+��6�.m���1�΅.�g3ZB�ek�5W�e��G���;_��8W�w��fDJT�к�&O�8�:�������P�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcNQv�GL�r����$lIdM�rv�BE��j�%@1��
_�0�[X�b\g�=�7�B�����&�\�e��n��*��.��P�&�}���ġ��,�4��[P�:ޑ�������1;[lz]G�ؒݷ��2Y�>�ԫ5�Y�w��2l��*��l���-f�8�[GB�S�j"Y�lK���;�>�k0�l��M���3�t���.˩�Y�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���X`
�e����1�:�Ω��x[,�Ns��{0��d#�t�  ",�V��o5]�Q;�im��ȍry��	w¹��<d���<
DN��$wq����+W���F�^�Y�7#�xI���E�����o)�]rH����8���f��9
�@�g47vΫ<�6�Q=h�5,Wlr�r%)cA�&�C�/�h��=;�_�8V��F�x)3پ������ׄ���MK�L�P�i2s�4<��!I��5��4]�폮h;e��w�5�ϟv�BA�IH���O,8(�6k�4d�Lt�2�t�U젩`#�4>?� �1Y��
�iC�&8�,��Q�L�������!�`�(i33��(b�W���5�.SƏw0�����98[Ɯ��X)�:O̐�V2XUt�{#	�x�=�tneX /*;63��dn��AmOeTky�q�\E��0</���/�u�[-�c]^�\�6m��G2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h���#}�Σ�f^ 
u2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�*���j��jR�o+ͦ��t������ׄ�:�CTt �\ ��q<qs�B�ӵǶ�	��l�N[�-e	�z�2������A��<��T0���S=�Z���6h�����s��Q��sr �����c���#R|��\�ݔړ��0������Ѿ��/@�qiQM��*���(%��}kutC������i{�W�G��!?�d���&�C#/<���q��3�*�M}x�C���Q�$�SE��'HY-m�@8��/=�e���-ņ`���"�R�7h�,b0V�u�Q�ݚ�Н��5���=\�B�wj$g8!�w� wk���,���9^-����y�,@���k���x�8�D"�����ׄ�R�
qtC�NI�Q4p�/Cj���C�1m�'*Gʯ7Պq�Y�.��x���"x�ś��5j�g��$P�M	�D�$ȨQ�?�Q,\ͨ܉p����O,8�ݚ�Н�h�'f R>N0Θ��ݚ�Н�Gظ0����t�%�Z?��<�ry^�%��C����\P�ʊQ�����J`�wӨj]h�vYv�������q��@����Mh?V��j�c�;J�*%n�+�uB;y��"Sek���6j�"Hs���%ˡ��V,b;�:��,����*���*-�,���O�]���N�����?�d���&�'3x)'�V�m7n,�
��W�.��A$�P������5d�������y�(����<m�r$ɓǃl[�Ƶ�1tSjv�?V��j�c3R�d�ܦdN�<@Iv��nt=:��:5A��p*qA����6\�4�@�� �-j�1tSjv��H�����}.z)yG��Hb� h�ҩ�?V��j�c3R�d�ܦ)�vL�����]W&fĉ>99��A0ok��$f��_Ub��7��G_��$�)�vxI��S�ud��E�9K��;_��8W�w��fD|]η����Αo��p2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc9Y���&���'܍|Cy���QJ�wk����\����|ݔ�3�(n�'�(�S��)��R�^Ƒ��;��|BEΟ��
�U�a�(��^GѬ�_���t�T��?E-h��`f���sC>��ӚH�RtV�^�'ž1�|�'����u��r��q�\E��04>^!b!4b�z'hۉ)��d�7�qĹ߆�p�h��d��JXl'�T��~��Uг�|<!�`�(i3��Nh�=f[���������<�.�����8��GM��-����!�`�(i3�v�Wס���G�K$x/��&���PC-��i0Q�͹�Ɩ,�b�R؅�!�`�(i3q�\E��0����G�t���m�� �ݪ���CyW�f�tR�wX��!�`�(i3��Ě�����}Dq�f��3��C���H�� �YߥթD�[*�Bi�v�V���;AD�e�{�W!�`�(i32+5�"�����-P��F����~�;2V-W��	c@�^ k�R�e�0���m�e#e>�=�^݊<���He�ylB��-t���m�� �ݪ�򈟕��+�v�7��]�ݚ�Н�3��0����g����F����~�;2V-W��	c@�^ k�R�e�0���m�e#e>�=�^݊����xQ�e�ylB��-t���m�� �ݪ�򈟕��+�v��t���?�� h�ҩ�!�`�(i3�lTN��I���q�}���{BO���5�%]���a(􆿳����^��!�`�(i3��jVѭ@!�`�(i3u?�:�H�jsrCm�k�J��6�d�t��w��X�'����u��r��!�`�(i3q�\E��0��@Z���rs�i�}�O��LTSG��ʎ�=U9��R�^Ƒ�Ӆ��I�ѪtR�^Ƒ�ӆ�v�9��!�`�(i3�����!�`�(i3�wӨj]h�(%����Z鎬�������(���/%Z�ڄ^1��#ƌ/B�ݪ��2�r5�����jV�{+�fbmDF�!�`�(i3���%>�rGO�D mWN!�`�(i3��Ě�����}Dq�f�HN��R��bP�63Z�tHN��R��bP�63Z�t��Ě����E�i�m}6߸��S�Ȍ o�n�J-�ƪe�0c�)�Ul����,�ǰ	r�R��Z����i�|7��_	�s�t�{���6������]'m���G�K$xE�p4rqG7]u��
�3�R�^Ƒ��;��|BEΟ��
�U�a�(��$��,Ix�6�o8:4�I���c�90B3v�A����èV\���F�`yx�>�+X�M?��y�!�`�(i3e�v��ҵl�{_8�Y��=�}�Vݨ��}Dq�f�����g�Z��3��a���!@�f")u��r��pT/�GS��%�����d��-��![L��^C�+a��o���H�RtV�^q�\E��0��@Z���rs�i�@24b��H�[���wkL�1p/-��G�<6�U����z~)���	6�
�:qEp�;�P�t�5fĉ>99��A0ok�׹�3��܌o��oŵE=��X�z��V��	��y�߬9�6ש`/V`L�v*2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc� ���j���Gɾ>�z����5Y��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�Y�Eat2�\��n�q�����"?��A$�P������5d��n4s1��7�癆cgQw�c4~Nr_�mS8<�n��!�3�
䖬n���/ ���we��0�U+�qbp@���{$@d9mh��n�tr�yÊ��_
�u}%GP����ZLN�	��� [-�9����G�^��D��!��"� +}0�ʂ�j�Ï��	�l�lM�3 H�RtV�^e<�Ia��la��o���H�RtV�^�wg�]��l�
@\�nQ�rV��q�t7��-����!�`�(i3�d�@���GU�lP4��/����*Q!�`�(i31���~�>=���#䖬n��؂�nF���<�W�.�P�	��
�Q�}HN��R��bP�63Z�t�G:w���he���!�T�1tSjv��>=���#��he�վɢ���he�U10���i!�`�(i31���~�>=���#��he�վɢ�F}���V6M��C��]��ġ��,���t+X�}��NۥUn��g��� �:5A��p$f��_Ub�F�S�1 ����F��O�}�	76�&�� Ӗ�t$�)�vx�J	���/a���Q=	+�{�*��{�ՖR���D�8�����t�T��?E-h��`f���sd=��¾ȼ\���F�`yx�>�+X�M?��yЃt����}����˃�I/ ���we��0�U+�qbp@��t����}�H_��#�Ր��V��e��0�U+�qbp@��t����}�H_��#�������i�e��0�U+�qbp@��t����}�H_��#�՚`��n����{_8�Y��=�}�Vݨ!��"� +}0�ʂ�j�Ï��	�l�lM�3 H�RtV�^e<�Ia��la��o���H�RtV�^Us��K���(yJ+��ʤ����3�W���b�0�T9��JG��NۥUn�+
�Tn@H�oi���:�l�^���;�jmT�#�>k�N��^��hJL��;���N0�!5R�u��r��;�jmT�#�����3�Ⱥ;
J��0�=<MW�-}�	mp5���%�+� h�ҩΪ���l���oi���:��*�·Op�r~�h��ݚ�Н���w�w:�!�`�(i3T9��JG��Bf����{_8�Y��=�}�Vݨ��}Dq�f�HN��R��bP�63Z�tHN��R��bP�63Z�t�Zj���
�d�@���G����B� �b��!�`�(i3�D���s����NۥUn��5��\���� h�ҩΪ���l���oi���:?�Bo���],��%s��'��_sN�">�������Ra])n#���r�����t����}�H_��#���վɢ�F}���V6��%��@qf���-A�¤�x.�Knqrh#��Y�
9mh��n$��k��3��,H/�����%>�rGO�D mWN���%>�rGO�D mWNHN��R��bP�63Z�t�5ߧE4��Fr��jϤ�Lǀ�r4��3m��Jw��3�+=�4o���+��+}�K=���e���Օ��qvdЧ^{�jM|�"D5�O�%E#P��=m緒1d�;q3�)�U��)���Y;e�iK!���d.O.C��|#HK��A(�c���_G��Hb� h�ҩΟ/��mS%y�W�CbE�{_8�Y��=�}�Vݨ��}Dq�f�	�)��&ghRV��RK7͍��|��W&":�;b�-�2�k+Q�h'�Ȝx�5W ��̫(� h�ҩζ
�t��T&���LQ�/81tSjv��B�'��a�S���%��������f��1.X!�`�(i3;d��'�XƤ5_���H(�T�O��{Tɀ�"'��&އ�[t�Y81�d�@���G�X���.��ġ��,H�Ћ�r�H�RtV�^;�jmT�#�YN
��)e���^b�~H����8�O�5���1tSjv�!�`�(i3�/��mS%�r\���%����g\>������
�:qEp'{w#/ B!�`�(i3	�)��&gha�E�Rq���my$�N��o�/���;!�`�(i3$f��_Ub�F�S�1 �fĉ>99��A0ok��fĉ>99��A0ok��$f��_Ub��7��G_��$�)�vxK���q
�&�lV*�]�aT��3G?�d���&���#��� �Rɫ�%�'�M��+��+}�K=���e���Օ��qvdЧ^{�jmWᅫw�5�O�%E#P	�)��&gh���(A�,"�(-w��N|;��|Bʦ?�H#F`�� �R�!�Fr忒@2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcۖh��)������E��㕷�f�Ux�_����+�b��T�Q5�r#�.�O 2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 �3 �����|��sQ�G�=�_�7V�o��_�Rv�䩲$��8��I�:Fa�7���z��O�|��/7*f'�|��bs��2[�a��o���H�RtV�^ϟ��7�4ÿ����Ԃ�nF���<�W�.�P�	��
�Q�}����g�Z��3��a���!@�f")u��r��܌;���'����u��r���Zj���
],��%s��ԏ ���ԭ�m��3��p���H���6Sa쎑t2�������50f
V��.ᬵy���Ÿ�`u�1tSjv�V�Ո��+5�4��c{�"�S��+�ϸ�i���U������՝� s�#���k$ ,��G��zł)w����ۥ�Y�mK7͍��|��W&":�ݚ�Н����F��O��;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6�������ł)w�����Al+�HB�����������mA�ѕf�f�_T:5�����2������}W`�J$˄���Z�׭ �k�3���u`�`�A ���\��o��_�Rv�䩲$��GQЌJ
��`���φ��<�6��ڱI�̘'np>�#�=�|#HK��A(�c���_G��Hb� h�ҩ�9�{�Jj3Ř�z��l �vPu06��K7͍��|��W&":�;b�-�2�k+Q�h'�Ȝx�5W ��̫(� h�ҩζ
�t��T&���LQ�/81tSjv�V�Ո��+5�4��c��W����W�/�#+*f|��sQ�G���+����rV���qޤos�em��ܑ��y���8���/�DY�7f�P:��z��l J	ibP�v
�:qEp�;�P�t�5fĉ>99��A0ok�׹���C���N�ky�A�掲t m^1r����,�ǰV6f����np>�#�=���-Q�OP���N��-��f���]_q�g�]@n_���?3Cy����]E;��|B����UrV���qޤ%�n#� �nF����bS��jarV���qޤܡ��F؝=��/z*x�n;��|Bs�'��OWnp>�#�=��Al+�H������B��/�����x��+�]'\gWg��	�Z�kfc�_	�Ƽ��S�J\7N2��j������mA�7�癆cgQw�c4~Nr_�mS8<�n���*y}ep8@)y@dl�SB%��I97��EN�h�h�u+��.ᬵy���ܝi���ؼ
���$����G��s��c�,��G��zB��/�����I(����K7͍��|��W&":����@|����^a�nu4Bޗ��jw�	���|#HK��=�O�-v�*_�mS8<�n�ݚ�Н�`)[�-hnhG�W�W�/�#+*fG9�:Q����t[�L�a\Y����+���LQ���"X��[��Q[R�7;�jmT�#~��F�����������yN��7��aq����i��oZ O\������U�._�nQ�rV��q�t7�l��8����aGl��Z����pG�p�P>M_���u��r��;�jmT�#`)[�-hn���+}ȵ�v��ONH!�`�(i3����ҧG9�:Q��� ɦ���AԢ�a\�Zx�.����#��o�TX5Ȭ7�j�W����^��D�Ϝ�}Dq�f��	��x��ݚ�Н�,��G��zB��/������R�s=Tu��H���9�-�a��W|!�`�(i3��Ě�����}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���ء�I��߸��S�ȌM��:�3��H���9�4���qB�Kj2�K����S�p�$@PJ+5����E�EG9�:Q���OLF+Q�>	#4�a��?b�@</�P����B��/�����>���Si9�i���>6�b NK�+���w� �~�^h�	�i^䖬n���n��y��a3}PR�]C$�.9�?	���58���d�@���G^?������X��O���r����!�`�(i3!�`�(i3����}>Y�&�-���k%�B��;���N���%�K�W/S��8(�E���Kt�emW��EG��-WBgW�6�h�g+�{�*,���H�z��ݠ�s����J��ͻ����8��Օ��qvdЧ^{�jmWᅫw�5�O�%E#P/Q]=��7�k]m��&k@C�Ɨ0z�cULj� 1�B��/����9-��g���t�
�:�WdM4@�r)1;�Os�rs�i��5O
T���ihc�ؓ;)Ve��˅�D�����R�`�|��K�z���k��$a(􆿳�3�m�
2]�����,�ǰ	M,��rER��p12���v1a{J�Զ �3 �����}c��ko#1^���E��'Z*)�?�R��nj��P_Q����t�h��W+��W�����"�>�3�eZ~��!���c�A�L'��B9[��EF�*���]�!��	Ǹ�y85���Ü�ۯm&����T��V��l/�#>6�b N>�3�eZ~��!���c�A�L'��B9[�o6Z^p�'���Xw�j�7��>6�b NK�+���w�(�)��c1�a-���7a
��r��L;Л����:<��j�.�g3Zv���� �_a���zz�2[QvA��q�q�ʩ)!��w������"��d���m��+�Z����y�{voPYӖt�iZ]XF�hx��G��N����p$��<
DN͗&8�,���o�|CZ�k]m��aFC��)k|p��z~r�X�<\�!�`�(i3�����
L�c�n�R�V�E�-�9����b���4��)+�[Z����&�+x��z�@CP&Aq�K�^��Q��G�S>\.�!::tm�0�i.�9�O�G?X2�K��2WI'�=��y0��s���4@Q�/���hy�NzK�}TR��b=���|��p��PIQ#�C,0�?����6[��u�9k�\,���m�
��,! �@��&}��{��Wӏ�c�ۡ�����*�v={k�h�+d�/Y�Z-u�e�8�ʫ�	�ϝ�YC�!��w��>6�b N�d���m��+�Z����y�{voPYӖt�iZ]XF�hx��G��N����p$��<
DN͗&8�,��@x��r�k]m��aFC��)k|p��z~r�X�<\�!�`�(i3�����
L�c�n�R�V�E�-�9����b���4��)+�[Z����&�+x��z�@CP&Aq�K�^��Q��G�S>\.�!::tm�0�i.�9�O�G?X2�K��2WI'�=��y0��s���4@Q�/���hy�NzK�}TR��b=���|��p��PIQ#�C,0�?����6[��u�9k�\,���m�
��,! �@��&}��{��W��Y#ѥh���*�v={k�h�+d�/Y�Z-uihc�ؓ;)	�ϝ�YC���*�)|/P2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcN%ڤ L���V��m[=��slc�)��3%�!Bd�&��p6(�*2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hW����Ga=]� X�Mgw�� gWVbT+踫g(�r�x�y�Zgl�k�����թ��H�V�n8�A�A�/�����y���|����4�[)�j����0��/�����T�
jl��.�.�g3Z�)V��B�1/������0�JB�� S�H͞ {�회�h�#5tNx�j�r�|2;$�JأͽgF"?nQ�rV��q�t7;��|B��� OD�C�x!�H���J��Ӊq��?Q�^�^E4+у��b�Bϱ����(�犽{Tɀ���S�<Ԣ��Oh��*��ġ��,���~����݁.�q�0��E|�,!|�α+N��	�Ȓ{A�dha#4\�0l�@��[����F}���V6JB�8^���m��3��p���H�����5{��&��.ᬵy���Ht�
�IZ�	|��9n���㬺$� %7䨅.�g3Z�)V��B�1/�����o�����;�|v�~�ٰ�Ř�hZ��~vV�V��j�3���xP^C�쌓�����&Y������ܤ�o�u�/����5X)m��p��I�K�#:��A$�P������5d��n4s1�U��B��-� �ѕC?"����z:fh͘�.�(�����xjzӝ���I(͂��-�����G�dE�h�k]m��F���d H��(ә��nF���<�W�.�P�	��
�Q�}W����G�iA'R�	��ೈ}�Ί$ԯ*�$)�'DV���b�z'hۉ)��d�7�q��k��^�1��dc�@c�����h��-�����s�Yls��8��GM��-������.J7h��C�x!�H���J��Ӊ}b��
��^�h۾�(�b�'Beͧ��&�~Lsf�e�}s�P�g�7�M^���H�L!�`�(i3�Ɔ �����O�����C�1�r5��(ә������D�v1a{J���ǔ���ǚ�F�d�c׮�1r���✯}Dq�f��5ߧE4��HN��R���ء�I��߸��S�Ȍzsلx1=�I(/2]�;�6*���'�
G/������Z� ��(H������D�v1a{J��;�6*��{%т�Zܑ��],��%s��tl��a�{q�����i���A�r�r+��½v1a{J��F��`�/�����sc�̆�!Y�X��9K��{%т�Zܑ��],��%s��y+��rf�s݁.�q�0��E|�,��	�Y2���Gg�&��,�0chC+��T�����D3���t�  ",�V��o5]�Q;�im��ȍry��	�
�I�>y!�`�(i3��i�\�{q����W�Ty��5��){�Ysy�t��P$u��&8�,�oa�}��p�-�o%�݃��x���Ԓ��t�2~?�������g�����t��:ҹ���7��I������-5Ԥ0Qo�n<�!s
9��
ss2����
)\Y�����'u���ɿJ�ҧ{�x����y�mZH֫&��5�q	�gh�䊉�䞘gx�n�W�����v;�k�@d���t��˳3[�u8�k/�z�xEQ���*[UxG�y��j��k
e�3+{�i�m�T�੉��%>�rG��M����{����"q�\E��0D������'���Xw�j�7���Ɔ ���9/�^Â?V��j�c�;J�*%n��Ɔ ���	�ϝ�YC�����%�!���Gg�&�B�~�aV~����E�+��@-�-'͏�������L��Hl��R�7h�,b0V�u�Qׇӭ�Ѿ
�I�>y!�`�(i3��i�\�{q����W�Ty��5���Fz��gCu(o?C!�`�(i3y�Z�;���>0�1ۍ�h �=��oٷU�b5�Όú}�ᛑ_��Ϩ�v1a{J��K�5OoL��C,l��e���z����M���ՊG*�؍��@1z�+J���5���Adu�5k
��F���U�hgh�䊉��	��J�6p�N��2�Q����:KG$��:�e�h�Ϧ^c!�6 �ef�v4=��/����t�$o'�Y��
�iCTl����
����P��0�&�ͭ�U젩`#���ٻk���ɕ�eY�����w6��&3+�-?V��j�c�
���!8Z鎬�������(���'�jh�,�cЉ�M����ve}(q�\E��0�sr���0/������K{��!ݏ�\�/\h2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!D� �B���9�V��r%֌�R����/7�o�H���7ӘK�!���{"?��	`��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�A��K��g��	���Ĝ��FKE|�q@C�x�>���� ܷ^.�c=��?�d���&�E���7-K|���|��йX#��S״$(�>g��������T�B�X
��=�_�7V�o��_�Rv�䩲$��8��I�:Fa�7���z��O�|��/7*f'�|��bs��2[�a��o���H�RtV�^)���A7�{�"�S�)P<�ܓ�Y�̢k���F�KD�Vr[/}>5��0�B� �b���H�����Yu�������&GV�Ո���VU[���I�)�ݳ��Y�Y`$�E�.1p�Y,CC�|^��V�Ո���VU[����� Vה�NEP�B�UB�I'?��t�Y|c��i��VU[����� Vה�NEP�B�UB�I'9gUS����-U �sȸ�"rR�Y�Y`$�E�4�B��AeO@�s��M��NEP�B�����n��}Dq�f��5ߧE4��HN��R���ء�I��߸��S�ȌM��:�3��NEP�B��Al+�H+*��xf�kUx���6�|����C�X�ҥՕ������}>p~z�r,؛��ap~z�r,k�@�&��T:5�����2������}
���!ꭶ��yN��7��aq��G�n���t�;���NI	��y7DT?�R��n}�����Hو����w/,�L�溥����v�8:ۛ@W:���#���F�P#�PC� l���E[J��:�������Н���˟��J5������I�?g�f&:��r-,>F�|��zʎ����%kR��������֢&@��&��x��&^�B�wj$g�X;p`��R<�����á�~O�,���9^-���.��֞�������i�-�;8|,����(��g.Cf���ϟ
B� �r�_�B&��p��ѿ)�L&�Fڱ���E�-�o%�烒�]������B��/Nߜ�*�l8�b(������l__��S1�c���Q��ǺΕR��ӟ-��G����JVW{�-v���m��3��p���H������7Pr��ġ��,Md*�;���D�&��� �4V�H�%p"��RR,���D�#��-�Vjo���po�h0�h�#"
s���
|�1�0j�K�^����\_9ͫ��Q������(���^�k��,�:�N�*�x3Lv	̅���X;p`�(�����֭�h��O5�tx\s�l.�	�C�
�:qEp��:��Zg�Hn7�(��wӨj]h�vYv���A�J�e�!�c�A�L'c�����O�D���|0f�?ǉ�=D�wP�/�w���bc��U�d�#�b�gD�XU���;_��8W�w��fD)IA����Cj����tLR�8ae�3J������ �a���GE�9TK��f�l0 ��J��9j.�l>'�o��&L�/<�t��Cn��P)��	�+�`g�]@n_���?3".3�]�N�L�溥����v�8:ۛ@W:���#���F��*{�욋�Օ��qvdЧ^{�j)�]�T��z�**ߜ�*�l8�b(������l__��E� )�&,�W�8"M�5�O�%E#Pڗ����7�9TK��̷_��yC��S8�vV�y��F�k]m����/z*x�n;��|BA��h�v������jֈ�U�d�#�bj�	17/+*��xf�kUx���6`�������X�ҥՕ������}>p~z�r,؛��ap~z�r,k�@�&��T:5�����2������})��uX�<��n쯎+�ܼ�P���(�K�g���yN��7��aq��G�n���t�;���NI	��y7DT?�R��n}�����Hو����w/,�L�溥����v�8:ۛ@W:���#���F�P#�PC� l���E[J��:�������Н���˟���p�;v�[�I�?g�f&:��r-,>F�|��zʎ����%kR��������֢&@��&��x��&^�B�wj$g�X;p`��R<�����á�~O�,���9^-���.��֞�������i�-�;8|,����(��g.Cf���ϟ
B� �r�_�B&��p��ѿ)�L&�Fڱ���E�-�o%�烒�]���f&m��K�hvl��9�h �=�'��L	�ߜ�*�l8�b(������l__��S1�c���Q��ǺΕR��ӟ-��G����JVW{�-v���m��3��p���H������7Pr��ġ��,�}Of��l���8��T�h���}둮j\����C$L$E�͆عE���ؼ(�K�^��Q��G�S>\.�!::tm�0�i.�9gh�䊉�䞘gx�n�W�����v����?�dv��oTN֢&@��&�_F�k-��苇��Fe#OOJd֯��|��p��PIQ#�C,0�?��ʉ��%>�rG��M����{����"�2��}��CϾH�)�]�!��	Ǹ�y85��J���K�+���w��@IAE�?V��j�c�;J�*%n�fePh����(.�G�k)���/z*q+6j�"HsF�prB/ˬ8��� �r-��M���>oKk�����jֈ�U�d�#�b��i0c���y>'MM귈nIg�R�5��/dV�ļަ��P���]6����(����c�n�R�HM���#g�`Bu�������}>p~z�r,�+�/��f���-A�¤�x.�Knq���;W��ZLN�	���M�X�FG�p�P�➁q��H�g 6ͥk�0�=<MW�-}�	mp,��_А#�<om��������oK?�d���&���>�9�=U�d�#�b�Dǁ��m�Y�{'%s��jb�ܳ�/�����b>I�WkxaT��3G?�d���&��!�k��w��=b��u�_3GH�F��7�Ͻ�{��w���Vڐ��$���юD���%�d����6����7}Wo�ָJ�}��;Nj����tLl�������'HY-��
�C��9��ϥ/5�����6��������֢&@��&����$G⃍�������������;^�6#9��u��n�k|p��z~r�X�<\�!�`�(i3*bL�(Rp~z�r,��Q�b��3�����}>p~z�r,um��x��m��3��p���H����Q#�?���;���Nå�a1��Y~�y�����[�5��H�o;<�6�Q=�	���c���KT
;��b�^"Bɨ �����V��m5Y)14 (�C0��٢�[.\�G]}�$C��� л�t�|̸9�73A}p��)�D�&��� �4V�H�%p"��RR,���D�#��-�Vgh�䊉��	��J�6p�N��2��,Wc��I�W�"�Ů7�6��,�ݜt��ϑ_�������� "5�]3Lv	̅���X;p`�(�������0�&�ͭ�U젩`#�4>?� �1%��C����\P�ʊQ:��IK��<��_(x��`g�%Y��̗0z�cUL#������b�'BeWh4:z�]MD�wP�/�w���bc������"d����.���k�y��t�+E���Q0�?mq94,�����5x�	~��TvukUx���6$E�?4\6B�@o��[^�}� u��O���#Q���< F��x�l��1:�N�*�x:��+���������i��@�����[�x�X���+���LQ�f�?ǉ�=�gCu(o?C!�`�(i3�m2��W�����}>p~z�r,E(7j�������}>p~z�r,���)�b�2������}w⵾k���yN��7��aq��hx��t�#���F�`�ã��Օ��qvdЧ^{�jb&P�"NE�<�6�Q=�	���c���KT
;��b�^"Bɨ �����V��m5Y)14 (�C0��٢�[.\�G]}�$C��� л�t�|̸9�73A}p��)�D�&��� �4V�H�%p"��RR,���D�#��-�Vgh�䊉��	��J�6p�N��2��,Wc��I�W�"�Ů7�6��,�ݜt��ϑ_�������� "5�]3Lv	̅���X;p`�(�������0�&�ͭ�U젩`#�4>?� �1%��C����\P�ʊQ:��IK��<��_(x��`g�%Y��̗0z�cUL#������b�'BeC���YXA�2��}���zgm##����Н���A�Y��|Dvܔ!�p�F�`n��i������+Z}͐�	}�@�r�<Uee�N�����$��̼�K���Z�׭ �k�3I$T�w�����+!�/}�u�F8O*�E`��f�A���yN��7��aq��hx��t�#���FӪ�c�g<;��|B�V���pu����p�5�"��[�B xh`�@�7�^E4+у��b�Bϱ�]h�(NAP/i�\	t�R��-�g� �GR��shbvk~�#x�l7�l�r�#���F��|}�&��3���.1t΀�+I@Lv�@[�JJ1��P�M��j�)6)-
3���WS=+E�
*��H+2siŞ�W�%3AԢ�a\�h�_e�8�4sg��ǎ�*��Zۉ�L�溥����v�8:hJ�tV�nQ�rV~��s�N�$²�ؗ$_Krt��qc�~�`롎q�C�r�X8g��mT�Of���-A�¤�x.�Knq��H�����ġ��,a��bt�eC�����m�������y	����F��،!|�α+s���s�֩h6$A����U��)���Y;e�iK!���d.[�����(����<m���"sS<�0�zG�������&G!�`�(i3v���,Ͽ�2[QvA�ͧ��&�~L~l�d����!���c�A�L'W»��`�{B�P��w(�f�� l��}I�?d�G5V������yN��7��aq��͹��e�[�.ᬵy����{!�)X+J��a�_݄:�fnp7Syv�Jы�^�)w������e��)��{}��M�+�'�̗������*��fPP!�`�(i3RnQ���_A}c��ko#)Ӄ�X��~l�d����!���c�A�L'W»��`�{B�P��w(�f�� l��}I�?d�G5V������yN��7��aq��͹��e�[�.ᬵy����{!�)X+J��a����P�L�E��w*��@�1�˓:�B��>Pi(���B���Q��ǺΕR��ӟ-����q���Ĺ߆�p�h��d��JXl'�T��~��Uг�|<!�`�(i3܌;���d��-��!i��$>�cQ׆��p0�Ĝ(�IyI�1"��f�Q׆��p0�Ĝ(�IyI�(�����'����u��r��!�`�(i3J���ٯHb�v��ONH!�`�(i3m�����Gd��}U؄�k]m�����m;
h�����B]�Pd��}U؄�k]m�����m;
h���^/�M2!�`�(i3z��-��g���k$ ���y��lDR�6؄���c�ۡ��F</h,��.�W	̷_��yC��S8����2Ho��@��@R�^8�*w��T��v�9��!�`�(i3
������}Dq�f�;�jmT�#P"G�wk��g�e��C�b�g����P�|T
�ʪܟ��[�x�X���+���LQ��B� �b��!�`�(i3�H����AԢ�a\�ۯ���@Z�2[QvA�ͧ��&�~L��X��� ��Cѻ�~���e�)qP@L0��U���(�犽{Tɀ�$����J�	�LÆ��S1�c������b5�2<B�!yf�� l����jA��L�L�溥����v�8:hJ�tV�nQ�rV~��s�N�$²�ؗ$_�#,���R�u��r��!�`�(i3��k�C�-�<�ao����O����8Q������51�X�c�rs�i� S�xSVe8��/��u@hy�`�w��v1a{J��\>Pq������^�L��,H/��!�`�(i3�����!�`�(i3�q�9�ͭhy�`�w��v1a{J��\>Pq�������B]�PZ鎬�������(���Y�&�-�yr�/ӶWȶ���/�Z�k�ʆ-�(i�pY%���m��3��p���H����HRCJ��<om���o�p��F��0,5 .�U%{.�V#?p�&���A �80D� �Y�]��`�E(���B���Q��ǺΕR��ӟ-����q����!�`�(i3��Ě�����}Dq�f����%>�rGO�D mWN!�`�(i3�5ߧE4��!�`�(i3�5ߧE4�퉅�%>�rG߸��S�Ȍ�M5b�&:|����*دHN��R��?�d���&�/�M�í��{_xGSn�����z����b�p����ī�����bL�'���IX0F�MV�ҁGG`5:�����+�^n=\f�5>�������Vmm�TF-���?4���R;�|#HK��A(�c���_G��Hb� h�ҩ�%��C���Q׆��p0~�5�H5m�v�&�k���������|e"%��C���Q׆��p0~�5�H������I*�&�v��/��kOT��ɕ�eYl�x���
��e���F7�Gh���l��,+)P<�ܓ�Y��+�t2�����dz����NR�p��@���|2Z��|��� �ҋ�;��}Dq�f��L�����B��2�k1�h�H��*��;�Â���ESҩ/��kOT١w��zj�X�X�>M�a���;}`O�k�4�����ˈ��`�@�./��kOT١w��zj�X�X�񳱅���^����z�嫋�T����|e"*qA����6\�4�@�� �-j�1tSjv��H�����Yu�������&G!�`�(i3&aD�4�X�X�[RP� .��ɒ�F��kB�t�x���@~H��k]m�����G�5����@~H��k]m���@� �
,9*�����
�:qEpNh���W<˥�'ܤ",�X�G[���7���B�t�x���@~H��k]m��E7�y�PjNh���W<˥�'ܤ",��E� ����e���,o�ݚ�Н�%��C���Q׆��p0~�5�HRoP��e�*�&�v��v�A�
^^3�V�C��k�HvL)��E��PT�Q׆��p0�Ĝ(�IyI�1������w5���iѹ�+�t2�����dz����NR�p��@���|2Z��|�����:l��0�5G,��Gc#����a4����dz����NR�p������jp����a�)�1�׀�<�6�Q==z!
���-�F�i��|�Uk�rDp!!v*!���K�5OoL!���}/
;$�Z��"�Y�<�SЮ!�`�(i3�L�����B��2�k1�h�H��*��;�Â���ESҩq���3��`��R�`K��"���վc7t��B��2�k1�h�H��*L]�f��e��
&YY��!�`�(i3g�>x�����H��6��b�4ƭ,�t��2� �צ�L��^�뢗�˯��Wނo̒.�9�lA�J�����١w��zj�X�X�>M�a���;}`O�k�4�����ˈ��`�@�.R��ak����`T�ҩ�	r�s�"���A���3A�n�+�sQ}b`�����E���v�RK��h�~s�K���Q\� C&����q��Z���Y�eF@�Af8�ٕ��(�W%����`ɊP�oT�L�ݚ�Н�?�C�KQ]˥�'ܤ",��Gc#�����O8��vW���V�C��k��38�h�3&���JT��ݚ�Н����F��O��;b�-�2��;�P�t�5W?�;��Ɨy�"c�z�
7!dB�c���Dx<�f�8ݵn����`Q�����^��h6$A����U��)���Y;e�iK!���d.O.C�U��B��-� �ѕC?"p���h����1�sH�RtV�^�'ž1�|�'����u��r��N
������Y�U��3Y��P4 �<�5Ɂ7dN�<@Iv��nt=:��:5A��pG� �l
s�M��KJ#�	g�˿��ji����{_8�Y��=�}�Vݨ��}Dq�f��L���������h\�L�O�c���ESҩK7͍��|��W&":�ݚ�Н��V��G F��x�⢄1@aw5�=Â��'e��0�U+�qbp@�!�`�(i3o� c �R�%1���%��K��>Pn��>�my$�N��o�/���;�B�'��a�'�7��E*��0U8��v��*����x����E2b�z'hۉ)��d�7�qĘV�52SG�U��@atA�ᴽ����rv:��q9+t�}�ݚ�Н��V��G !]�~F��A�mi�K�7�����//�ƍ2���lę�k�C�-�<�ao��6���z�S�yC�wbN�dN�<@Iv��nt=:��:5A��p�e�<Q��Y#ѥhZiC�������;q�{_8�Y��=�}�Vݨ��}Dq�f�I&!y'}�}c��ko#ƌ0Q_,�I����~uK7͍��|��W&":�ݚ�Н�^)�G�B�+�WdM4@����[y�K�/ ���we��0�U+�qbp@�՝� s�#0�ʂ�j�Ï��	�l�lM�3 H�RtV�^܌;���d��-��!i��$>�cQ׆��p0~�5�H������I�I�߷�c/��-����!�`�(i3����6`X�/m>8Φ�ʽP�Rܷઍ����:~�Y����.��������h�4��=y����͘6��q��kUx���63��<�����ݚ�Н�G� �l
s�M��KJ#�	g�˿��ji����V��G �pȌ���]���E:�qL��n��p��b�Bϱ�fePh�����yf sg���}Dq�f�L��/\��=2���H��̣��O�˰�]q8k��.ͥ�H�RtV�^��.J7h����ly�P�r��n�Ŀh$�*�]�`�,\��ݝۺ���r��������]�Y�_�H��!�`�(i3�����!�`�(i3/w1z��ӊx�D�Re|����xت�����:~�Y���Wql����BM"���}Dq�f�HN��R��bP�63Z�t�V�52SG�U��@atA�ᴽ����rv:��
w�	������9�~�gz��8�,�@�VҒm�L��@�a��Hb�2�Ǐ��Pn<���@���(9[���G�������+��<�ao���#!��H�ȯղ!�`�(i3v���,Ͽ�2[QvA����[y�K�Q����!��Hb�2�Ǐ��Pn<��!�w(�y?fĉ>99��A0ok���H�����Yu���*Y��b"Wfי�b����{�6�o� c ��f� .):_�mS8<�n�ݚ�Н�t�R!ME��ߦ?�~F��C~/*�t�2�q㬑u����p�5�"��[�B���p�8����Q����.��$���g�e��t����3��v�9�ʘV�52SG�U��@at3Y��P4v��*�����*�R���Amr��8On9�*�����C.�u�X��I�ՠ�w�O�����|�D���H���~�����l���X�� QT��0+��?�DEu�>��-��4�1tSjv�!�`�(i3af��pD�Ї�6~��Ȕж�{�7�^E4+у��b�Bϱ�����ס�07Syv�Jы�^�)�:5A��p�Ra])n#���r������.J7h����ly�P�r��n�Ŀht�2�q㬑u����p��8��V\⯜�'�,LF!�w(�y?
�:qEp�;�P�t�5!�`�(i3�V��G !]�~F��A�mi�K�7�_�R��U��@atA�ᴽ�R܀{�!�`�(i3^)�G�B�+�WdM4@�%ρ��r�}6�/S� 8��/��u@�n�Jt�g�v1a{J����w �!�`�(i3I&!y'}�[��m�Uƌ0Q_,DE(_
/�n�Jt�g�v1a{J��A&��R�����%>�rGE�}�Wk�m�ڨ�hծHN��R��bP�63Z�t��ܐ�}Ď���!�+����=@�Hhg� آP��n~���=2���H��̣�� �<�5Ɂ7^���H> ���8ѳʳAM��KJ#�	g��7������Hb�2�Ǐ��Pn<����5��-�����dz����NR�p��@���|2Z��|���-��4�%m�Y$� 1Q#�6q�U��@atA�ᴽ�t�2�q㬑�M�{�|L��!ߩ��`4%�fZF�Gck��x������=l�H���3���� �����G��D�h��y@�Af8�ٕ��(�W�5���^�.I�����wl53�e�%^oe�Y���q��w�X�X�񳱅��5��]���h��N�M��z3:��K�z{�� ��C~/*��f� .):����6`X�/m>8Φ�ck��x�����ٷu�/��kOT�n���h�n�&Sq�a;Uйc�e�0�RAL�!hy�`�w��v1a{J��]%���0��8ѳʳA���9�~��� �������xNetҌ5`��K7͍��|��W&":��u[���ew���m����x��O rQ��qD���FD>�v��Pn<���S�׫�hc�!ߩ��`��0+��?l�/��X��MV�,oF*�L��!�`�(i3!�`�(i3!�`�(i3�q�]��~S��b�Bϱ��Y�X-�jjL�E��w*�8.����6_f.�}�ٷ/Tu����W`GU�!i&G�\��u���9�9��g"c{r�Va�irR��ak����`T1�h�H��*�������fF*�L��!�`�(i3!�`�(i3!�`�(i3k��_� ��(ӈ���l4Z�/��m�$����F�f�J��K��>P�a��]�/֢��s�Kȓ�FG���<���+tx�D�Re|����xؑ@�VҒm͏ڹ�)�u="��x8I�t�2�q㬑��&g�hh\�F�u������ހ�af��pD�Ї�6~��Ȕж�{�7���LM��Q�&�-�8Q�F���"�>mS@*�1�:�Ω�����|"�4ԲcZ7��n	l��Q;�im��ȍry��	:��+���������i�����+��cW���}���i����0���LO���){�Ysy�t��P$u��&8�,�V:i���ߜ�*�l8�b(��+�w]�B׿�ġ��,�b���30�D�&��� �4V�H�%p"��RR,���D�#��-�Vjo���po�h0�h�#"
s���
|�1�0j�K�^����\_9ͫ��Q������(���^�k��,�:�N�*�x3Lv	̅���X;p`�(�����֭�h��O5�tx\s�l.�	�C�
�:qEp��:��Zg�Hn7�(��wӨj]h�vYv���A�J�e�!�c�A�L'`���y��֢��s�Kȓ�FG���B7Ԅ��{k�h�+�0��NZ�Hb�2�Ǐ��t�搩�՚�(��ؾ#(�[�(D��_�W�F7�Gh딶�<?�3x�В&=�y�q}��2��*��t�iZ]XF�hx��G��!�`�(i3U��֜��3!�`�(i3X�PC!v�@[�JJ1��P�M��,���9^-���.��֞�������i�_o�dZ � �GR��shbvk~�#xǩ"�4s2nQ�rVA�H��%��SFU� �hΡKCh��(	�G��^����K�7����&Y��V�ǣ©��$��:�e�hfH'��!�i����VZDf�?ǉ�=�O�G?X2�K��2WI'�=��yp����nZ���t��˳3[�u8��M�g����H��bf�?ǉ�=̇i�d�?�4�0 L?�p���@Z�6[��u�9k�\,���m�
��,!q�\E��0D������'���Xw�j�7���ڹ�)�u="��x8IȂ}�5N@!�`�(i3@ E���߲	[F42�Y#ѥh���Ƭ��,��i�X�:D�o@~��=��X��/���Ȣy�!�3�4�f��<�ao����O�������R��j���C.�u�X��I�ՠ�w�O���/+�>�m!QFc��ݍ��FD>�v�t*�����b�氦�=��X��/{A�dha#4�8�e
��'�i�*ڶ�UKs,��l�?�C�g_3GH�F��Ll��_�]���LM��Q�&�-�8�<�ao��8C��D9�C3x�В&=�y�q}��2��*��t�iZ]XF�hx��G��!�`�(i3U��֜��3!�`�(i3X�PC!v�@[�JJ1��P�M��,���9^-���.��֞�������i�4��%�;��g��cH�wA�?�W��7E��n���8��T�h���}둮j\����C$L$E�͆عE���ؼ(�K�^��Q��G�S>\.�!::tm�0�i.�9gh�䊉�䞘gx�n�W�����v����?�dv��oTN֢&@��&�_F�k-��苇��Fe#OOJd֯��|��p��PIQ#�C,0�?��ʉ��%>�rG��M����{����"�2��}��CϾH�)v���,Ͽ�2[QvA����D/@�2��}���zgm##�v���,Ͽ�2[QvA�gN|���!|Z���wj��89����Y#ѥhB�@o��[^�}� u��O���#Q�4ك��	ቢ��S���� "5�]�D:���@���k��!�`�(i3Y��B��7Syv�Jы�^�)f�?ǉ�=�����ݱ���������%'`�T:5�����2������}�k�+9=��@1z�+J���5���Adu�5k
��Fɴ|�O�j�gh�䊉��	��J�6p�N��2��,Wc��I$��:�e�h�Ϧ^c!�6 �ef�&�2�������ȍry��	Y��
�iCTl�������l6���0�&�ͭ�U젩`#�4>?� �1��ɕ�eY�����w6YmC,igu?V��j�c�
���!8�@��A���k]m���
�s�?V��j�c�;J�*%n��@��A���k]m����"����8�*i�$�HV��	��y ��f"���py�+��;����w�R���y����C������R첖쬽oj�΁!�Fr忒@2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�ų�Mƶ��^�
Q����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�#�"-�vz!�`�(i3B�t�x��')6��;��W�����/
���aː���>#��0����3��N��x]-�
M�<vW�9�+��NЏ�s_(1��P�=���6�ĢZO�}�1U��VP�CXm������>?p�8Q"yM��V!�D�WaU�	�D�6I^��V���u��[�,���E%4��l���M���R��ӟ-�F���ˏ��Z�כ��c0zQu�<����i"��@#('�cH1��<9Oy��]#�0D�	�I���_
�u�_C�7�2������}0n�V2���]#��t�ѕ1��ŦL�ݚ�Н�!�`�(i3!�`�(i3پ[���-��Z?�6j�"HsضZ�i\�ώ ���]q<���}c��?:ͪ�'g�Dw[���/=��Y��Բ�@cD�����L�#}�{���j�3�����M�ë�fBz��|2���U�����vl�-p���Og����n�貶|?��R����w�����@-p�h_�=i�/����#���K��>�;�0�j�?���+���͵�p�����g�����q(��չ}/������Z����
���\hW� *� �}�����1mS�Q��v��$#d�bu�r<���}c�»�<+h�Ԁ�~˼��H����8����F)�~��[t�Y813bQ=�3�� �֤D�A�m\�����Z�כ��c0zQu�<����i"��@#('�cH1��<9Oy��]#�0D�	�I���_
�u�_C�7�2������},��������yb52�_�8g��.ᬵy�� �a~�"�;Q١Ӿ�$w���	�e���0��Qܓ'{w#/ B!�`�(i3!�`�(i3!�`�(i3��%>%��w�R���y�sL]~цt�U(i��[�,��(��F[U��=��YV�g��L�*� )�\�~xyf�-�b�{'{O��c_`J?�R��nj��P_Q�[i_1|`�S޲�U2+q,� L���?�q0-p;��|B$  ��$,K�9+�/���p��\��be�����E8R�c4!`���U�._����P�|T�ݩ^�H(�BM�ܤm|��R�TE7SmQ١Ӿ�$w���	�e���0��Qܓ'{w#/ B!�`�(i3!�`�(i3!�`�(i3��%>%��w�R���y�sL]~цt�U(i��[�,��ᥨ����a)��K�Nl�x����b�'Be��
����Ѳh��N�M��G��-y�� ����i9v�A=K�����_
�u�}���:D�_�k�Æ��%N��� �"�W�A�&hH\m�:�5P Hߜ�*�l8�b(������l__�c�9ʼ��$����Fp7�D�_�k��HM���#g[|��;�ċ�lʥ��|�]v�A�9I��@������Z>��~��l��"�
k��x̥�0�L�p~z�r,�%⠩��!�`�(i3!�`�(i3!�`�(i3?Q�@X>#�[}[���Q׆��p0�Ĝ(�IyI �q�T�<�C,�#1��<9Oy��]#�YUw�d��F}���V6������X�hvl��9�h �=�{UY�Z�[2�h �=�'��L	�ߜ�*�l8�b(������l__��S1�c���Q��ǺΕR��ӟ-�G1������j~�]�������:�.�{4\����^��.��8?�o[L��h �=�����=��/R�c4!`�d>�c�n��N.�6��9��t�i.�#�),s=�����}>p~z�r,�q1�G��o>0�1ۍ�h �=�)��=���!�`�(i3!�`�(i3!�`�(i3?Q�@X>#�[}[���Q׆��p0�Ĝ(�IyI�h#"�.^����p
v1��<9Oy��]#�YUw�d��F}���V6������X�hvl��9�h �=�{UY�Z�[2�h �=����y|���D�_�k�W�A�&hH\�LZ:�\�Ԋ�{Tɀ�$����nQ�rV~��s�N�h�5,Wlr�r%)cA�F��=��g�]@n_���?3ֳ���[HDȚ��wz;�|�����I�HM���#g��I�mV�Z9I��@������Z>��~��l������IV���@�\#��hvl��9�h �=���_��')�c�n�RÆ��%N��ݚ�Н�!�`�(i3!�`�(i3!�`�(i3}Y;�jn��~v�9p��0�5G,��Gc#�����0o�;�6�E�u�N����dz����NR�p�'q�-��nEg�N>Z��^�T��렾�������S�L�0�5G,��Gc#�����0Ö�΄�*�E�u�N����dz����NR�p�'q�-��nEg�N>Zϕ��<w렾�������r=8 ��FD>�v�ހ�mcW�ɓ�>0j�oc.�d�Y��~SC�	��%�Y)���N�N<҃&��;��|BG�r
�ɞV�C��k����?dq���z����7�Ia���^���H> �0c���cͧD��_�W�.��;�#��&�qҸ�2Mz`��B鼙y��ԭ�m��3��p���H������7Pr��ġ��,u��|zO�	��%�Y)���N�N�ƥ�FJ��?.��N[j��/z*q+6j�"HsӅ�X��^�Y#ѥh�g8V#��4֡\�`!|��.I�ܨ�@��A��2��� �s[�v՝"[�ya�i��{�7{�2z����!Cu�>(���] 9��)�
p�"��d���!iZ�,��#�2
��e�������m[�LEE�S��-��h���d�0���.�g3Zꢯ�wv��n�Jt�g���E�*��p�O2!?����^�� �|ֳ��V2-+;X���1�#��d_!�`�(i3� ��U�_:�[�qaV�7���a{����U�._����P�|TDqId�ja�<om����F6̜�����a{��d>�c�n��N.�6�����k$ !�`�(i3?Q�@X>#��ŕpO"��d�jO)īIX0F�MV�ҁGG%4vkz����`���φ��<�6��9;��ˉy��>>��A(�c���_G��Hb� h�ҩηxmQ,ۘSk���������|e"ʬw�S����F�n�8���[{/;k+Q�h'�Ȝx�5W ��̫(� h�ҩ�y�}�6f&rG��Hb� h�ҩΌr���h�0�I����~u#� �,W��	��uc���q�D��1���~���Z�@���v�;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6��9;��ˉH�ٌCx�`	HX'�}'����g��cH�wA�?ܵ��� �?�d���&��]�o��A����\��]8��	���#�z��%]'\gWg��	�Z�kfc?�#	*]]�iI9�o«IX0F�M��ŊPTWo9���b��|2\���F�`yx�>�+X�M?��y�!�`�(i3z�
1���;��nF���<�W�.�P�	��
�Q�}�k��^�1��dc�@c�����h��-����;�jmT�#�,l����M?��y�!�`�(i3���J�^�G�yd����f�m7�IB�>9gUS����a$�/�4�	��E${5j=�����%>�rGO�D mWNHN��R��bP�63Z�t��ܐ�}ī��K��M�ZP�����Fz��Ԥܑ�9�ڮW;��|BC�5,e�������'y��$�t�Щ��I��gs7ߐ)�~ң>0�1ۍ�h �=�,�W�8"M�5�O�%E#P���J�^�Gs��>H�,b�z'hۉ)�4�	��������w�R���y��0�J����e���?ͧc� x��p\�>�7���o��_�Rv�䩲$��8��I�:Fa�7������A����ᳮ�T�7�癆cgQw�c4~Nr_�mS8<�nx��7��G$�ء�!�`�(i3!�`�(i3!�`�(i3��$�\%e��}Dq�f�v�A�
^^3�V�C��k��Q4� 
!�`�(i3n��>�my$�N��o�/���;��ɕ�eYl�x����b�'Ben2WȔ�h!�`�(i3x����E2b�z'hۉ)��d�7�q��6[��u����@~H��k]m��n�_��-��!�`�(i3E�g�������(ӈ���m�r����t�R!ME�D��_�W�.��;�#��&�qҸ�]b ��^E4+у��b�Bϱ��L�溥����v�8:ۛ@W:���#���F�Q+o�>u����p�����+X��FJ���-],��%s�����F<j��.#�#�-�p�@�Af8�ٕ��(�W�!Ċ&���X�G[�,<���g�F}���V6��%��@qf���-A�¤�x.�Knq���;W��ZLN�	�褩�23p\� C&����q��Z���2%�ɛ'�F7�Gh�8�n�"X��:5A��pu����p�����+X��FJ���-3L�*}F�J�a$�Y dN�<@Iv��nt=:��:5A��pu����p�����+X��FJ���-��]�q�J�a$�Y dN�<@Iv��nt=:��:5A��pZ�,��#�2
��e�������m[�X���2:#J�a$�Y dN�<@Iv��nt=:�$r�t�}ik+Q�h'�Ȝx�5W ��̫(� h�ҩ�y�}�6f&rG��Hb� h�ҩ�t�R!ME�!�`�(i3!�`�(i3׾ŞWsuz�6�<������NM�����ɕ�eYl�x����b�'Be�&�����S&aD�4�X�X�>c�.A�(��cS�c�X�X�>c�.A�ݵ�Q�n��T�\ �͉ק��l����@~H��k]m����s�>���ݚ�Н�&aD�4�X�X�>c�.A��`���TNh���W<˥�'ܤ",��E� ��"U�7s,�/Tu�����_&������@��9gUS����a$�/v�A�
^^3�V�C��k�HvL)���D��� �!�`�(i3v�A�
^^3�V�C��k�HvL)���t��GU�Wfי�b��}!D̅��t/)����(��cS�c�X�X�>c�.A�L]�f��e���"X��[b�&�,���Nh���W<˥�'ܤ",�����D�-��1�K�!���aR�!�`�(i3q���3��`��R�`��ƍ ��s�!ǵ�N����dz����NR�p������jpR�n�G-������+X��FJ���-6�5Y�S;a(􆿳��3��TY�@�Af8�ٕ��(�W�!Ċ&��V+���]7�wtMM�0�5G,��Gc#%@Ԫ┇	��*��\� C&����q��Z���Y�eF@�Af8�ٕ��(�W%����`ܑ��y���8���/�>�h��fLD��_�W�.��;�#�E���_	��}Dq�f�dl��[�����{�6�*F=ॵ��@x8��vW���V�C��k����?dq���z����7�P'9�V�˥�'ܤ",����^�� �YW;C�͈H�=��
ڨg��U-�e�%���/�X�X�>M�a���;}`O�kй�Z�>���;b�-�2��;�P�t�5�H�����Yu���*Y��b"Wfי�b��}!D̅����<!GO#(��cS�c�X�X�>c�.A�x���0�������Oݥ��{)�h �=�$��bY\���ZAL�:y�g��K��7�I�$Q�ϐ �S���pj; �B�o�+�m
Og:Ba=�u��Y'G�vw�B��qbb��fddf�ݲ�UC֬g'�J|���������k{s�^,ysA�U�y��6��3fU����O���X#��cA;�jmT�#u����p�����+X��FJ���-],��%s��?,[�����v��ONH!�`�(i3�L�����B��2�k1�h�H��*F7	G�<�*�P�ߚ�6���}�%DܭD��_�W�.��;�#��&�qҸ�]b ���G�x )HN��R��bP�63Z�t��Ě�����}Dq�f�e<�Ia��lb~*��s�&aD�4�X�X�>c�.A��w�`�f�(���@~H��k]m��+�<;"��}�mH��q�=��Cn��P)�`�m���wa��o���<N��ig�+�?c2JCI��i�pk�<cm^�Y�F���_|@k�q��Z��}��oC�H�"�]陒(Ѡ;�n-i�\�*�ߣ3� >/��7�I�$Q��w��b���u��"����ٰ�Ř�hX8�P���C�X�T�b\��ݚ�Н��ج�B��\� C&����q��Z���2%�ɛ'�F7�Gh���Z��� h�ҩ�7�wtMM�0�5G,��Gc#�����0o� c ��Dǁ��m�@�Af8�ٕ��(�W�!Ċ&���X�G[�����K
�:qEp�;�P�t�5fĉ>99��A0ok�����F��O�\E�W��4bƗy�"c���c5�^�H"X�0��n���l�IX0F�MV�ҁGG%4vkz����`���φ��<�6�Q١Ӿ�$	��1�h\���F�`yx�>�+X�M?��y�Bz�;{/�>��]#�y�W�CbE�{_8�Y��=�}�Vݨ��}Dq�f�Y�)�}��EXs70��nF���<�W�.�P�	��
�Q�}����g�Z��3��a���!@�f")u��r��܌;���'����u��r��a�F�������Y���D��3��b�]결���:$�O���jF�ཕu�_�mS8<�n�ݚ�Н� �#0xg�`�I��Wz}�ἱc��-).^QQ�b��~$�
�:qEp�;�P�t�5����l��~��?�kv��.V��:��������kB�����X!o%�ſ����O?���/�4�j�`�;���N����?�p1tSjv������$�D厺��+�̟�14�����{��O?��ʔ��,Vr՝� s�#���k$ ����������zՠ�����˦G�K7͍��|��W&":�ݚ�Н����F��O��;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6�Q١Ӿ�$�C���j��A�����P�U��)���Y;e�iK!���d.���+�^n=\f�5>����Db^<�..�4���x�H@�[xjzӝ���I(͂��-����>�Q�c6���*(H=�ƍ2���l�����g�Z��3��a���!@�f")u��r��܌;���'����u��r��>�Q�c6�~nS��\z-+;X���W���b�0���Ě����E�i�m}6O�D mWN��ܐ�}�~(�����Z�@���v�j��A��4�	��������A$�P������5d��n4s1�U��B��-ն'�U;|�u}D��Ǫ2�q�m�bs��2[�a��o���H�RtV�^�4�	��3|v��Eb�z'hۉ)��d�7�q��k��^�1��dc�@c�����h��-�����s�Yls��8��GM��-����;�jmT�#~��F�����������yN��7��aq����i��oZ O\������U�._�nQ�rVj����vy�B� �b��!�`�(i32VP��Ѣ��P@JɈ.���3R��6 y2��R�	��x��ݚ�Н�EOJ�uxm�7d��2�4.K7͍��|��W&":�ݚ�Н����F��O��;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6��R�7ʌ�J;\�6�{�ѵ1�c�{���w�|@C����8��Օ��qvdЧ^{�jmWᅫw�5�O�%E#P��=m緒X�X�pF�{_8�Y��=�}�VݨaT��3G?�d���&����*�����n��e�����u��&Z5˞�� �#1@h�5,Wlr�r%)cA��z>9�R��d���!itB"o
�B7Y'��k���=R��Ԗ�A$�P������5d�cp6Dq��;���EWr���e�T�5���u�L�xZ��j�
�iB{�Z�_���}�\���0�=<MW�-}�	mp�?IK��y�8���/�l|�*"k���(ӈ���m�r�����$�Qu�������l3��K�y��Fp����f���,(���B���Q��ǺΕR��ӟ-�F`���G���Cҷ��eV����(K7͍��|��W&":cp6Dq��;���EWr�kv޶Gl��d˵T�d�٣��c�A�L')�_��rT�`��9d�R�e�0���e A7YzE!�`�(i3l|�*"k���(ӈ���m�r�������+�^n=\f�5>����Db^<�..�4���x�H@�[\���F�`yx�>�+X�M?��y�!�`�(i3���e�T�5���u�L��ˇ�h��<�W�.�P�	��
�Q�}%Q�[�J3��K�u��>���e��0�U+�qbp@�!�`�(i3�kv޶Gl��d˵T�ˇ�h��<�W�.�P�	��
�Q�}�k��^�1��dc�@c�����h��-����;�jmT�#�,l����M?��y�!�`�(i3��=m緒�`�	�l.�;wjN�rs�i�E�8�w���P�nq�S�p%�t;�{�B�'��a���p��b��]c�)�#y�D�5�S�`�	�O`�� \)�H��������P#o�]�ʄ���e�������aGl��xF�oͧ�ߜ�*�l8�b(��MdGN���!�`�(i3V�ؗ�X`u!/��"��E����8U��@�fћ���Fa>t!�`�(i3�d������)���܇�b~*��s�͝������XƤ5_���H(�T�O��{Tɀ�"'��&އ��-/a8!�`�(i3M*KJJ�[�4br��l|�*"k���(ӈ���m�r����!�`�(i3�I��� g3��K�ޅ7�=w�'�̗����S]�_�_��u��r��!�`�(i3	�)��&gh?d��ǧ�C�|J3J�n �v>������
�:qEp'{w#/ B!�`�(i3	�)��&gh?d��ǧdN�<@Iv��nt=:��:5A��p
�:qEp�;�P�t�5!�`�(i3���F��O��ݚ�Н����F��O��;b�-�2��;�P�t�5W?�;�끤g��ޏ�S�G��T8�q���uҽw�R���y����<�..�4��M���|c��'��*��I.��^�