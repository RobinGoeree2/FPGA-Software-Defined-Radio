��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���G�H�ƻ	�"�iQ�����3�7Q��㼫F|�ݽ0��@h ���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�S�T�;Ϗk[�^��_���Q� ���6��H4ي��2_)��:B!�b�ؐ:�{T�{df�r�<�XD�* O�:��׶��{�*Z���H��ea�8���*���g S��/P�p��]��;�I�����)O��Ξ4�"�\�� ���K�O�{��
2�D�� ���Jc\֣�I��B���t��|U|�/֚m� �+d��.8%D.��n�P��<2�q�U��k�8u[\E���@N1�w�0XL����[fe�Hs��9lSUQ�S��)���2Ee�Y�R2
�I.��	���
����k�������0�?�}4��ѕ�������U��=>bMab�	;4��G����a�����(�I�?g�f�L#����2=�l����3�����U���T�����\�4�sc�[�.����(�Y���mG�z���_15~n� L������ѥ�Q�hʢ!�5�bAg�
d�m���i�h}�a�mC�0�Yf�Y�F.�"�K����	x]�m�Je{q����3U�Ƭ8�5����B�3ʦU��&}Xa���qd��.ݫ�hv��m�!=�y����h�}T��nJ8��>��PY������kGQ��2��2�~�MUs ���7a�N^��)Y.��]�ߏ��P�umSe��S�7�׫X@Sϛh^�X/���H�3�g��Yr
� �AH�T�t��3��'�Wا[�[?���̾J KNW>�F@�4%��Њהt�#��Zhǀ�Һ�3{����V���	x]�����O�Я�mڍ'T����X��Hߵg�:�%�+T%2q򋙔�M-US-�8<�n�У�Ǝ!�ѠV�>!�/�7��u���nEA~1�a���;t��⫓���RL�a)3���ʉ����H7�Q?�"�B��@�$�;�7C��H���j�v�?�r	⚎���k�8���҆�|n����vJ�^�R�!�"s̊#�}��uJ�Й�m�BdP*4�h־�-9�,ڸ@9����c�.[K��mN,����0j Oag�ì���Tl��!���<< �sN۪�c�	u�~Rp�,k���%k�&ָ��sE��D�őⴔIꈸV�MT7xB2I�d�HnULkIh��:h
�[ϸ��W�A��S;CM���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcz��9�L����WS��]$�Q�L��S����E@��~���($�J.���
�=W�֯��i@F�5�=h�GD�#�̔"v��ƒ)?˳R����.��ѬL�1m��+Y#_WӢۉ���2=�l�����4�c��ҁ�o���h�k2�$�����(����5�2���[@%����nEA� ��]���\"�&@�4'���Xwߍ���y�CV�6IWJE�r���秹��ч���2eI�gxBo�A;h�F�`�"Q���]�!��s�XZ8E@�KXϔ�×��̙̳=-� �`#��.X���*"v%)�(��(����������A�=���ѝa�l߱���Қp%�;��0����GI$��ǂcY�~�s<��MR6�q����*�JvW(�%��b����i�Ӛ��F�)[ Z|X��Z�H�(�*�b�βł1Y�ΊS&��$шe1Y�ΊS&������'l���u66�v��G���`���o���"��y��� ����;*��k��J���\��[CK�VsC�~��~���+4������f�^i�h�];�����X���P\�q[�7�����a�"e͉�Xk_�0��'nU�óM�˄No�M����f�g�n�(�r`M�5�:v�9/��=��K�(�+k�y�_%��5�J*�Rs�0_��T��·_����J�	�LÆ����Us����M��_(����@1Y�ΊS&Q$n�ti�`������3�V2����"u��֦5d[RM��A���D]�$���k�1 �O�o������*���ɪ�{�e,I�!���7�mdy�-�AG���^`	��x���AC'[U�7�tW-�J4p'�>��\��:��Z鎬�������(���w�?�b�>��]�!���٥���E[U�7�tW-�J4p'�>��\��:��AԢ�a\�w�?�b�>��]�!��u���Ʊ���T��xdE���ƪϤ�Yk"1/���%	v3�t�  ",�!�=��F���"�|�E+��T����oGo�Z�J��ݪ�"�却G��B)�6��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�pv��[�\�)�A��m�aOLyb�7�a�`�2G%�/��Z>L}x��=��f0���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc\�BDL���iM0�3y��#Q���Q�q��o
�X���C�~��~�Ln��S�W�ѐw���5u�0�yo�_���
.����Ď�rȫ�S ��Sup�xg쬉� }�ֱ�q������m�q�.4g$�co��=��ەI7յ[+8�Ǎ^�~�篯����hV$��-�����$�[��= -|�GP�ݚ�Н�
ҭ�3���#���1���b����@�Y~�`���Y-]�\^M�Ɣ�	��x��ݚ�Н�
ҭ�3���#���1���b����@�Y~�`���Y-]���v�9����Ě���!��"� +}���k$ ���n����-�����y��j��k\y[P޽��5 cd���%��E�/�xA���%0[-��&J��;b�-�2�'{w#/ BƸv��*Qx�!F�;^/K�2�+����e
,�p8�4��|r$J�-��^$f��_Ub��7��G_���;�P�t�5�37y�����:�3��s���EU1��?�}����0�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������P���2�z�I0���ԏc�r�(���7L��1�6`3bQ=�3��>�Dj�OgW���y�k�m2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ����"��y��� ����;*��k��J���\Ol����֑1Y�ΊS&�<�ɰ]�+��׌#��M'��P+V�_������o@i�1�P\�q[�7�����a�"e͉�Xk����0��hC$?���;���EWrf�Nd+l�Yҽ֗�1#��Z�����f���T,m����i�Ӛ��F�)[ Z|X��ٖ���g�OcH��9d���aX���$�Qu�&�<��G�!�`�(i37w|s���0�$i��kq?H^��2踫g(�r�N�ǁ�f�T��p_U
#yO�E���%�;���EWr�L�����!�`�(i3�b9���1]�?��� ��b�FP&��"��IJ�N�Q9�����-�)����=��ەI7յ[+8�Ǎ^�~�篯����hV$��-������"�=�X|�\dG��&(i�/B�\3���l�c1���~��DFTޱ}���0|Q�>8�ހ�$f��_Ub����b���잸��u��r��>���(���;*��k��� ��y���Y-]�[�Q0�M�1���~_'R�4���%�3�F�������78�4��|r?\�z?Xk�:䩒=]'5�����}Y��	}�@�r�<Uee�N������*��vbsQ?M8�f2ݜ�
N#�0���:s����"��IJ�N�Q9���2��n�v��/��@���#��M&s��"��IJ�N�Q9������وt����jVѭ@�y��j��kj�����N��L����͜�}Dq�f��5ߧE4��L�{	����Wma9h8wc������5���!�w(�y?�?�JY�)�Y`��jD4�7�癆cg���&Bzv��`f�(��H�RtV�^RD�+����N�ǁ�f�T��p_U
#��ʟ�1G@<�6�Q=ٌ�{m�tOIkV�g�ػF:7��*W�;֒	��x�(�6k�4d����Fi��I��RhF���9���x��
&\C��J_�0����O��Ě������������0u�\k|RSm�y��c!�Fr忒@2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc>sh�ڌ6�ve���'�=�9���bg2r0b�wa�!��@o����8����`4�+��+ER��{ia,���ߡ�c �ج�γI�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc.�
͹U���|K�{ߝ�Fc��B�I%ji�7��
#>:��� �rmd�&l�����i�I��M�3q��=$���A���ۖ?3�'����1Y�ΊS&nQ�rV�kV�џ�}$|~ïSup�xg쬉� }�A�%��fOX��8�r�;T3���/�"[Ʈ��JHn��z�F�x�aK�k��GZ>.�004@�k8���F�5/K �*jE|�ڴ�>��Xӌ��=)֞�)56s@��t�N�}�`�k��?Ŗ��R�A�%��fOX]a��1qh_�n�To�[�C��-��JHn��z�Lqܳ<��J*�Rs�0��(o <[J�	�LÆ�ѯ�x��yŮ���z��!z2}s�Uʚ7�ܩ�.fOe	Ln��S�W�"Lq�q/��Q��ǺΕE4���0Q��J���6�,A)�ؚ�����
��\�H��/Sg�w��'op�[�d�3���`�kq͠|�zDN�-�!I��'���N�"9���b�=����r{d��JHn��z��c�Bo��F:����Į��KH ��ߞD�ǒ�J���6�.X��;;"����v������*�%� �2S��(_�<��=k�Rm���Yci��zW�F:����Į��KH ����멋��I))����A�m�(��ʢ
w��]��0�ȍ�x�>c��w��'o�Q�kŕ��Q�Ӹ$P���F�׼K�3
�v�v-}�	mp̮�%I�����0i��Y��f������&J�b, ӫ/��m�B�K��1Ҹ�]��0�ȍ�x�>c��w��'o�<���q��q+����>(\�H��/Sg�w��'o�6���OB\�Ns&x������F�׼K�3
�v�v-}�	mpl�!����_�n�To�[�C��-��ɨ]^(���Ѹ���_�j�`���: ��ao.\C�k���uf|ò���
��_������B�K��1��n�da�ۣqM��X�~ ӫ/��m�D�K�h�x#�L_ѭ�Q�#3�d^�ϓ��ͬz�Ť��!4�%�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ�oZ�o�S��	p���DUeH��lW"`oG&2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc\�BDL�t�� ���OgۈPML�����"{�B���}$|~Ð�BY
���wb�S��V��^��\i�ֱ�q������m�q�k�v_Q�(��Қp%�0�ΩyO^~�R���ce���n��8&���I���|I���:�Ϊ���L�8ɵ��i7N�_�M�3|r (���B����}�-�f ���:=��1���h�E)�.�2u�ɯ/wI���?����}�	76�&�R�Q���~��p���웂���a�"<b��5^,��*V�m��'��3�V2���i=�d����s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�i/F@���V.F����R��kBޫKp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hN>�4�
���y[6���ڀN�&jl�o2C�g�kgw�"��I��R� V�pFr����A"�U���w�c*����W"��ό���.�d=��¾ȼƸv��*Qxm�QA�Q* 5�����}Y�]��h@�YyZ��}�Q?M8�f2$ Hl�]��u3�0~͗��3��}�	76�&�R�V�"�0ɶ37y�����:��Y�g�f��߼
�dUY��~�6� ��5}�Y7s�9���o��S8��@糺뾃7܌:����3Eֱ�q������m�q�>1�Pq�@\w��0]���8-|�Dp��xs�S�)P<�ܓ�Y��=�g���>��8��-�Ϡ���:=
ҭ�3���VFc�B:�pO���w�_fHN��R��Gu�"�0�R�@�6�֐����o����(��e鎃9���1�L�]�b�֘m��+��$|��;D���J7"(�=3Ի9|