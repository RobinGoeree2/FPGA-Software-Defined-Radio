��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���G�H�ƻ	�"�iQ�����3�7Q��㼫F|�ݽ0��@h ���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω������?9X�1�Z�U���T��ײ2��>���^k�/7�?1�(�c��ly[�$D֍C95^T��6\Xa��7��Į�N��=i�@x_\q[�@�0�I���j{�N<��;��� B]�pE���	x]̃Dj#^Da����M���Af\O��x^Q\7�z����)�,�˛D��w���旴4�����<��a��rl�ʩ{�Bfळ��)���X�$� ���jǎX������n�q��}�p� �Ñ�]�*�p�㈍x�!����Y�f��a�Z��Vb$���N[E�=����tL��	Z�G�a}CK�fC���4�O�"�F�È���_�O��<$e|����w'��1�:�Ω������?9X�1�Z�U���T�����\�4�sP	�b\qB��������"^Y怄����v�~�MUs a"�x���2@�+���c�#s�0���!Z:���:r�a�u�����!�M��E%<�$�7.�/��aG�k�8���҆�|n���:�o�E��Uu-M�rt�d{��}lJ�Й�m��?�Vޱ������{����VjrHS�w�MH��j���r���+W��YJt�,�y"r� J&g~���c*& z�s�ђ�B�~f��0(�/��$ }2����T���Q���!i��ӯ�02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vce��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�׍E�+��
���*,f$�7Q0- ��Ck�fÜ�2/���}����сsU%���n��/���Û�E�tw:g?�y��h�I����uk1i�f1?���b1�F��,��n�2��C�`Qe�IC�_�\H�F?t�)�Y¹w�.� -��E�I�?g�f�Jm*)�m��+���%	v3�t�  ",����%H�$��ī�o��<�)�G!�u�����!�M��Evl3����SO,F=d9�[l�&��q�©���H��JnXeS5H�j.F�6�Z��'i��'p�@�I�?g�f��Qө}�i���W:SJr���S��:C�-�䉢��S��(�B4�rs�F�r�f�t?�1J&�|D�e�!��L�D��6S�]V�H7'�R�^Ƒ�ӥ�e%)>�Z��&��J��Vǃ���O�4ۤ�`�	��B�f�\�kA�/����<.+6J!�t���\�Ws��l=�L؅��FJ��G��k���؍��R��j�.(Wx*9��?xs���}�ڍ������5	��]�!��	Ǹ�y85��1}�\���;�¬pX��g��U-�e�,���6+�^�9.�JQ!�`�(i3��{l�f|��rs�i�� ��*b��0��E|�,�CyW�f�tR�wX�Ռꢤ�Og�?�e����]�!��	Ǹ�y85�����څ��;�¬pX��g��U-�e�,���6+��A�y�0� 7G#+�Ǘ0z�cULjaGkƊ~F˯�+)�"j���b7���Øf�XA���BU7Ê7�E�4'���Xw�_�!	�\�����5	��]�!����M[��Ǣۧ2���{�ҋX����>��l%i�-̇i�d�?���{l�f|�ό���.ӳ�
�	?�<7Ê7�E�4'���XwI<��f�@O�x�7���q�©�����<��������S��R�9��0�S�&�����"m�K7{�>P�2-i_���F�� �yz��$6ea�8��������?9�f�*ʝ��R;�{m�B��Ҝ��a�N�}��t_���Յ;��n�a�x�a(􆿳��Ak�y�y/��=��K��]z�Sk����+��_�F�����CY���<�;�L���9��Xv7�j�i���TR�^Ƒ�ӽ�}^v��Z鎬�������(���`$�P.eE���lC��U�T�\ ��i3�|)sՀή.mH^�+��@}�M�`t�A~h}Nw��諚��y�[��0���߫�]�!��	Ǹ�y85��1}�\���;�¬pX��g��U-�e,%�0g����Ed��>�^);�OA�uW7s�9���o��S8�J�]=��R�^Ƒ����"X��[��Q[R�7����n9읃g9l���z��Q]� _�rs�i�jf� l�Ǜ������CyW�f�tR�wX��}�
�?����om)��%��(��+'���Xw�j�7��ct�:��RE��W��_�ړ8���/��O���O��ْ5
�8��S��?�F��SO�P��P����&��B�"p�l~V��o5]��lO ܅d�� л�E��QvfZ!4Я\�rƛ�}���1�)�c��!�`�(i3�E����F�Z�>)�ώ�~+�ݗ����>[H��_0Vձ!�`�(i3,ԯ���gn��Ab�%^��}Dq�f����gRI/)�ak�m6�E����F�Z�>)�����˟y���!s�;�Rn\�_c����L�{���D	��U�l>o��|��P�^/�h���/�dSƏw0���wN��0]fH��>d]=]A��O�T=�4e=��-Y�VN�=�ԕd�tuшb��jߺ��0�5tU���+�J��U<o^.K�}/��<Ӭ��|#HK��@=���b��0�5tUзq8�Ј)w�<�_N`E�cvR+��}Dq�f���R��V���X�&�E����F���8�TP��@E�`�8���&��Ŷ;���I�PD�na"�,�>E��4];ˍH����TI��Ԫ,щ�"��<H��(����O�c����L�{jݭ�F���p� o��]��hy�/B/���^!�������>�s�/���U<o^.K�}qW8+����8���&�qr�^*4y-X��;^�8�1-i4];ˍH��E�(��n6�Ѯ� л�U��v��;fZ!4Я\�rƛ�}��k�-i�9~�!�`�(i3!�`�(i3,ԯ���gn��Ab�%^��}Dq�f��N�v�1��B�r��!�`�(i3,ԯ���gn��Ab�%^��}Dq�f����gRI/,�Xʚ@h!�`�(i3,ԯ���gn�J����� ��}Dq�f�{p�R�I8$vVqYY!�`�(i3���D	��U�l>o��|���JLm|��������A?Љ'�-{<qH�~�!�`�(i37�ܥ��2���kܪ���*�LNm�d�tu���ād�,��x��B5�!�`�(i3x�]�V����:L���2*Q=F��:УWKŃS:H��+܆"BT�(���B�r��зq8�Ј)w�<�_N`E�cvR+��}Dq�f�{p�R�I8��a�=L!�`�(i3���D	��U�l>o��|���bǬ�='�u�uX]�Rn\�_�B�r��"�,�>E��4];ˍH��\B�����g�q~[{Q��`�)J*;�p�aٓ�v1a{J�*�8#�������8�TPm=_g}b��t�֚S��~r�S\w���!�`�(i3зq8�Ј)w�<�_N��M��+?���C&���t� ��Oz!�
�W@!�`�(i3���+�J��U<o^.K�}/��<Ӭ�/�"����J^L��z!�
�W@!�`�(i37�ܥ��2�`e7��9��×�>��|�\m���X����,�Xʚ@h�E����F���8�TP��@E�`�8���&��Ŷ;��z!�
�W@!�`�(i3=]A��O�T=�4e=��-Y�VN�=��7p�J��PWV����ftj5 8��!�`�(i3jݭ�F���p� o��]��hy�/B/���^!�������>,�Xʚ@hx�]�V���t���CՐ3��F<Y��j3��� Q�N��*���������c�] S�4];ˍH��E�(��<���A�� ;�Ӆ�&�`�����k@|�%5'��E����F���8�TP��]&�Hž_�FȘ�i��Nj�,�F�v��@���z\�m���Iϕ������z_۬=�!�`�(i3"�,�>E��4];ˍH�C#��N;F��D]�+�~���{/��I(�c?Hh�`K]!�`�(i3!�`�(i3!�`�(i3jݭ�F���,Y�y^:�3�y��j��k��V��e�LtW��e���d�tAAI�O����07�ܥ��2�k��`����VU��d�˰8���&�-�_��>H��n�-�!�`�(i3!�`�(i3���+�J��U<o^.K�}��HwL�X�|#HK��fu��n�!�`�(i3!�`�(i3!�`�(i3���D	��U�l>o��|���z>�n�S�|#HK��fu��n���H�1�� !�`�(i3!�`�(i3���D	��U�l>o��|���z>�n�S���*y}e��?=�2����o��!�`�(i3!�`�(i3,ԯ���gn�J����� ��}Dq�f���R~�e��ד*�h��F�v�C!�`�(i3=]A��O�T=�4e=��-������yM�8���&�9��^K��[N���b�����sd�!�`�(i3���+�J��U<o^.K�},ufOX�mCž_�FȤo�f�Ԝ��MU�@!~�X����Ѵ���X:��+�
H��m��E4];ˍH��1l��m�ئ��b�􏮚ǖ�!�����T"*�M��d��p∺V��܅���9��ȓM�Me����OA�,s>w��Bw�B�"p�l~/�"���꤭%�3��{�o��C!T*p�VU��J!�`�(i3!�`�(i3!�`�(i3"�,�>E���� &N��nF�d����
F�`�����1݁mP2<WV��
i�c�r�N>�X�5G�7Ê7�E�4'���Xw!�`�(i3!�`�(i3!�`�(i3!�`�(i3)��� ��1����_<X����"�����q��l0+���yn�����門�ҋX����Q��C� ��!�`�(i3!�`�(i3!�`�(i3k��j �%j!bM�9�&?�>�M�O�IQ���}t�{#	�x�u��߹c���o��C!T*Y�{'%s��F���u@����]�7�v�ԯ��Nb-�h�dN�<@Iv�,.9������:5A��p��1���P�Ivu.rg�q��l0q�\E��0���門�ҋX������S8�=	���/|2��#�	�T�\ ���KD��}[e��0�U�S{����<�6�Q=�qő��{XҹvXI)�vNd�)i�'�al��p�@��O���Z鎬�������(���pu�˂�tj{%��ߛ�8���/���}Dq�f�F�d����k�2��J>eR�<�V�Zt%��m&<�,0 ���Ţ�{l�f|��rs�i���YN���o#�_T��,0=]^	�&Z�n��[��{_8�Y���˂lq�㜯}Dq�f�F�d����4�������eR�<�V�ȓM�Me��aL�!��t�j�!󊾵�e�;Pq]g\ ���ǋҠ7�	�ߥ�H�^ /m�6���<�6�Q=���Ң�Q<�6�Q=	I%Mq��`Ҧ�׶!z1��,,ҹ�$�OD��G͘��P�!а��K��k-J����:M���FM�`;$�l���1��in�uM������A��[B�)�b!F��9�����Ïb�}������c�.D�#�ҒIs{�>Y��}�:_�_5:��(�I>�IP�b������:�kR�$fOyQ���؟�-�X��_��n��&�P��00�Ͷ\��[��=<�6�Q=�w�3����f
�@"��g�����Mgs�4�H�O��	�� ��Fw"�Ş|H��S��q<� �77AƐ^�8�s�٩�삢^��)('���Xw�����U���=����t�kD��*�ҋX����L$�����/���%��Y�i`YS����O0�P2<WV�����F�eO�V2y/��S:�cN���dt�{�Yi`YS����6+W��!�`�(i3!�`�(i3<�6�Q=�U�"���M]�B��5.��$�]��tK�"8���ɮ�� л�B)vظ�u�!�`�(i3!�`�(i3���y��lD�U&"���+c��k��Vj����C$��*V�ֆ�\��[��=��hy�xl��B �i<��z��}�<ͧ�:|�"��ӌ�r,�ttT𔛨Z��ΣS�)37J*u�,�JL���*��c�d}];�SSyZr@u!�0�"� ��w� 9_�똣w�ٽv�yq�`0�|(O��"��"�T�>�#�ҒIs{�D������:_�_5:��(�I>�IP�b�����LQo����������0��]㯟�Ķ��d����;���!�v{:��h�k-J����:M���FM�`;$�l���1��in���� zԻ�弳$_N� ���ui�X\�̈́nlH�I<�6�Q=���x��<�6�Q=	I%Mq��`Ҧ�׶!z1��,���F��qJ�?�̃�*�`��n�E�T����X�=���P�;�ȓM�Me���T��G���X��4tΘIy����ߗ��L1�%TԞ}�{J��n��&�P��k<kbm�t�vc;?N�ʡV�l�竷b��"&�=��(��Z鎬����Ĺ#{����}Dq�f���#:�LH�ҋX����L$�����/�����z|�\m���SLq�N���@��O���Z鎬����Ĺ#{����}Dq�f��5Nleo��ݑ���<��z��}�<ͧ�:|�>d�g�K��I(�c@� ��<��z��}�0z�cUL9kX����_G��?g��ORuD,0=]^	�&Z�n��[��{_8�Y���˂lq�㜯}Dq�f�F�d������~�~�8�1P��#K�SM0.�>k0��0ǽi�*��]�!��	Ǹ�y85��q幊s�?����H�c�B���)�g��U-�ee�@Rv����my$�N��;� ��b�� л�d�q=N$,����hQ���}VA�ڦ�c4�RP�m��q��ˑ��N��k�I#�\(z:�ĭ3S��n��@IE�U����S8�=	���/lg������T�\ �́��Wl� -��J�x"GeY𶣂���S.��TD���rs�i���YN���j[��v2ba(􆿳����r
��qő��{r��  <�!�d�<8�c{}�x���� ��6%j_�zl</�'.�w�4z9Z��E����F�_V�VG�88�;矷��N�����?�d���&����q��w);�OA�uW!�`�(i3!�`�(i3!�`�(i3!�`�(i3�s���6`� �3�<�G%�MP3$�x�Wt!�`�(i3!�`�(i3!�`�(i3J�a$�Y F�*3���6���Հ^����I!�`�(i3!�`�(i3!�`�(i3!�`�(i3A����2�2�h�8Vb5�J��>q�'�X�ǎs�&I/B�]���o��_�Rz���n H{y����i�q,?5qM�>Fr����7|)�`�H����Aj��t�35L��$
8��2�ֈe1tSjv�?V��j�c�[N�&ѐ!�`�(i3!�`�(i3!�`�(i3����;q�V.��(�t��5(kL����Ě����E�i�m}6߸��S�ȌM�>Fr���X�ǎs�Ӑg�(O�b��T�Q5!�`�(i3>�w��B]'\gWg�3[{���:յ[+8���,8?<�%�z�-uͺ�s�η3G��Hb� h�ҩ�{k�h�+��=C�u�!�`�(i3!�`�(i3!�`�(i3mQ��RA���oz�N��=y���ؔ���,�P�ԙ��i����I����l��jZ\C��>CM?��y�!�`�(i3d1E �s�)���Q���3[�u8��a�}�$�&�[.ǣoJ�ܯ	�J3�iU7��{���om)����5(kL��HN��R��bP�63Z�t��Ě����E�i�m}6߸��S�Ȍ��8�8!s��ڻC�i�;��|BK�B�<�t��I%U��_bM+���C����
&h���ٙ���O�Q���*��P�Vr���F�!��c���Y�҈�FQ��ݢt\�y~?��t�iZ]XF�hx��G��!�`�(i3D�c=p�^&�c��J"HƏ~g��ղT�D3H	�ݚ�Н����-��?s�_{X4u�`'s^?n�(�tc���u*_���X1'1[���A�|���$y̮�K��v ���X�u�Ӛ&&ĕ^$&B6�mC��[���ԗ��6%�a��x��&^&Y�o�wd��X;p`�ct�:��RE3z%�u�܆N����p$�Q����͗&8�,��w�Iſ�Κes��O!�`�(i3�nxL�J�J��2����^��9R�^Ƒ��f�?ǉ�=M7^��T�d��y��$wq�����0��E|�,
�e�~w�J3���;�_�������� "5�]��'T���+%�����-��i�m�T��!�`�(i3�v1a{J��H��S�A�J�e�!�c�A�L'1Ջ�=t[�}����SƏw0��;%.T-��3H����'���Xw�j�7���Պ�t$�;f�?ǉ�="]�ϓM��!�`�(i3>N0Θ��ݚ�Н��@����M>N0Θ��ݚ�Н�� 䉇o�M���w0�z�Gb��P�!�`�(i3B)vظ�u�M몴PBoT�ݚ�Н���O�q�̍!�`�(i37�_M��f�?ǉ�=����G!�`�(i3�d�)bU\����Vv�	�6���Ic����L�{�f%DR�*�!�`�(i3��/z*x�n;��|B��)���i����i,(��*>rc��08�����4C����#��̻�Yi#���!�`�(i3(h�+Z�RL;p�����@�ۻ����4%��0/�'�al��p���K酦z�Gb��P��O����Y��(�
t��Y�{'%s�Ǹ2����E�vwx�k�g��U-�eI?��b��C���/S�)37J*uG(�~ �,���cZ�����o��C!T*�q���U�<�F@"~�@� ��<��z��}�0z�cUL��Jv(K�V��c�4��s���o��x�8���/����\�����A���I��{l�f|��rs�i��s�٭�`�̳��i;��m�S��T�\ ����m0��~�bO\�Rэ�ҋX����7�8����u�c:ɶ��o��C!T*Y�{'%s�Ǹ2����E�vwx�k�g��U-�e��{����w5���ݗ��]����$)@���S��?�FH�$a��ma��bft������y�;���g����0ж�~a��bft��N���m��;���g����0ж�~KԂ��U=��5��L�����;�줦,���<C���O�G��o��s4k�r�j�b#[�o����x�&��'�|�7����s�ݺᣄ#��̳�y�5`P�~�s��hvo���$y̮�K��v �
VWk �0=�b ��"r1��?t7u�`'s^�`}��AyE=�b ��"r�?i���7�|s���q��W�qd�'��n�1��ņ�}h$�ɹ��I���x:����aR�!�`�(i3(T�流����>�SS�]n7A��^⠻rRV�������.�lz\�Q��?s�_{X4x�]�V�����TI���0D�Ub��g��~�4�"4D�/�k�_�|��|�7���@*p?{n��*�LNm�(�V*�u���ƸL��؅��FJ��o�C���j�R�s���-&J�ULnU�x�]�V�����n�l�z��q]4-�k���n��F[�e.VJHn��z�ʨ�lC!�i��}Gz���.��6ǿv�ɢ������=���a��z>�n�S�['Ȑ2��;�Q~���A�U� ���_Y�VN�=��i��}Gz�������vy�|�7���@*p?{n��*�LNm�|��yf{��������K�� ���i7�ܥ��2�/��:M/�CՐ3��F<@�Bcj;�J^��J�Y��h]^"���x�]�V���E�(�� �TYD���`
^8L���o��x�R5�A�yx�]�V���E�(�� �TYD���`
^8L���o���	L]q�x�]�V���E�(�� �TYD��BY��I��O�䓟�&ݏ��A�7�ܥ��2���C�0��(����і�Ʒ��u7btcǹ8ߗ:w��@!~�X�X�]�v��� л�ԭ:h%~k��u�������b,/^/��ux��:S?v!�`�(i3�E����F���8�TP--M�pu�����]��!�`�(i3�d=}b�TY���t�!�`�(i3!�`�(i3%Ah�%4
>��XP��ȆS�%������=�-�o�F[`3*�!!�`�(i3!�`�(i3!�`�(i3�b9���:&�>��s�� �5�v�^*?�z�̒�7�dz�H!�`�(i3!�`�(i3"�,�>E����\�v��_�R�G���Fz�Ͷ��>��9	�F(�Z~}�U��!�`�(i3зq8�Ј)w�<�_N��M��+?�^qk�d	��2Y��kک�)��j)yc�n�.�_�t����ˑ���M��iT1Η)say�s��l>o��|���&l@�[�ݸ�OK����DK7}!�`�(i3���4����4Ieŉh!�`�(i3!�`�(i3%Ah�%4
>��XP���{���r#�LN����p$`�̳��i;v�f7)�!�`�(i3!�`�(i3�b9����4�6�t�!�`�(i3CH�׳�B%