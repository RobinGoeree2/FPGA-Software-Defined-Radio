��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����⽸���D��6T�8�{N�/i�kf�!�6��̋"X��:�����\N(h�-����}!���1�����4�0���S��k��Xd�d���{�8�%���AHǚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>>�Htdʮz_�0�`��@�[D˂8��k�ľF�n�Ԥ��r�τ�u�&&����\l&�$������<H�����}�ƌRS>�(B-~�� ��ڣ�9#M��c��&��C:��pSv@1�{=\�4T�K�ݣƐGm������t�T]fē�����S��H/Am-
H3�6����	HK������%�0���&��D���tq3���Q�A5d��A_����2H3�5�J�K|&.>��ny�6�-�]&���t���g%�7��c��s�_�v6�/pY@�Sŭ�M*%�����q���8C�@0�o	��b!��$7*�a��,ƴ�Y:��q�%����
�6�E��(���Nyu�AȤ~�t%t:=�z)��0���w�Y���|�9���gJڝ� 5�T�sS��Q�mb��м����\zGd�:����Z�F�֐ru�������)��u����p�6*lً������aGC�E��;�*���M�h�k١���A�ȴk��3
�P0�R��#��o�-~R�|��k�*�`39�?��L8;4�g:�p~�u��O���Ťj8G+nut���T�Q �r$5b�n���-�n�h�
���^[GB���:;��E6ߎ���f
V}��K^q�K�<�9�prY�S�a�ċ�(@ok�2�Y:qIv���9��oAE2�qU�P�H�����Fyh��$OM%�zZ7�4�f���T1O�S֪�|ƶD΅}���D��^���<�m�'G�,�,o�X�tO��#���ɂ��şA��BA�r�	�g�B(Jz���m�ק����#��+t������S�7{��>� �/>ٜ��jL����T��̮- #��N_���"���+-�P�H�u���eލ����Ĵ���&:�N9����57��9^��~$i>a�!i ��#��C��AN��� "��ac>�"����MJ�D�E����};XN��_�(�+g2?�Z���$���H��}�x$�6�,��y��)
��kU�!E=%���!|����@�F�y��.�`>^��6���7*t���.�$f�F�}Y��DyP�
N��2�My�0�!��d����?aZF#��y�p ���o��Iߪ ����b� _��I��PA��2�������횐�q��J�x������KC�U %� ]U]W�G�f��h�u)u�!�ǣ�� z��=������O�����F֟��P@�\��ٜ,!�� 	���E\(PŅ4�F
,�>��ü�Ӭl��h��7�3�T��k�C ��8'H��J*Z	J3�>!�:\A*�/9m)n���ϋ���H��1�\c[Qa�F��
�#%q��{���m��Dtnv�b�(��P�,n8��͔pq6!O|�'������8unLUl�ѐ�̉��cB*�|��ђ�{}|�.T5���C�h.J��q��X��X�avGO�����	1���M��4�3?��o-S ��xmFܤRb*�e�����q,&c�yy�'�*70|��֜�V�=!lK�Rd��
-t����;��L�(�t�-�r���͊wE8�1� �@_�y�>�@����T`I,4R�o0�{U��L�8�\��Ua{����(17}7�Uc���]l��#�u�����Ż��ԡzuGo!0t{ד-�`�M�\<�^BW��Ǖ�����~��Q�}�nmX`�/,%�A����B�nњ$�?m{=�����%��<!��z��;{z����Ts�J$�g+	%�����~�����C�-���֢4x��;֌�
& � ��J�D6�'0;у�qM��ѕ~���:�lu���f�(+�ۍ״��t�:jᶞ�8|��c}0Jȁ5��%%�J#��C�R4�a�^���>QL�2|} S��e2E��Th��k�"��+����Ew��d�-���Qӱ@�b�?�w%Ӝc�5��^�/k,SZ�C�S"�h��<��\�)>$(���k2LsQ���]����/�
d�Tbؖ�7��*m���x��J�(���c�_��Z6��%�X�v~���p�ѐA>�L���МULy��/߬w�WJ��1K�[;�n|м���M�:cV:R@F�/fԛZQ4���;�!n���5���#댉�z�D�1{�\e%%�T�	}�t�wD�Z]|��?y���rU�*���l��LK�e�jJ���P�N��=I:�6��������s/5�~�J���%O��:n��j����(�ȕ��-��Oxʔ�/�e���rIa�ٛb��E ��+�_�\X%o�nB��燃�f뭈Ӏ<?���2F47�W^w^k�tW�筵��w�1 ��H�0��gt�[�S��i�4�,�Ϯ[��]�y�F�:����2L�F']��C����}�:�?�u`����_y��gf������v������=��X��|�XPlby��pJ�����+���Rx��n]�7��Jn'ɸ�}�U�?��D�2!�s�P��Az����[sR �;!��e�����Y�S΅$�X�0� {Ɯ ��ĿLRTc^�|�|�x��{|A4��i�X� �@��M�d�'Cw����	��+�~H�K!�bΏ���I���T�_�ٛ��RS�9C�Z�H�����������ے,nB�G��m]���&�SC�k+�E/�.�  ����x�w_�W��{�o�K�T�(�
���C�ġs$X�S���4�!������@��*��0���0X��F~�Ԗs��(�\1��-�ا���S=��U��l����f� AEή��7k��3�Ou5�Ё���_��y�|Y7za�.e��F��SʛL8� �41���B��/r�<c+��'�r.�[i)gX҅+�,`|uA���z�c��d'���w��������jY�e�c��礰��;�d�u�2/'�X�Y�N(خ�p5��dP���Xt�����'���~f�3�ӛ���}"ڇ:�Ǝ]��uc��m�c}0��%�$>I����g�J�k�S�RwS�t^H�"a�Cw�9ԙ�I�?��x�$�˚�lr/����,�� �eD���S)Wo*z���|��X�!Ƶ:���m�a���9^�,��]������	 �Zu1w�A���o���,�!ۯwx�@����Nk����Y�W�M�`��ͤ���C�R�#�j�t2�+�3�� :ҺU�,�I͢Q@�%�r�=��pZD+r�D���2*