��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����⽸���D��6T�8�{N�/i�kf�!�6��̋"X��:�����\N(h�-����}!���1�����4�0���S��k��Xd�d���{�8�%���AHǚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf^��$�i�g�Wɐ�)
�Ql�Y�+6�iѰ�^���d�u�.�Ye�ZG�$*�f�pM��Y���f<���YB�H6]��^�8�G{��:RjeQ��2
�ƣː��5JLO%/.�)����\�
,��YIw_�aJ�/��]b<Q�	{>�nP?/;Rqd�ӓ�Vn3~���Z������������J:��n��� ��j�=��8H��r�t��F2�t^t9��*�^R3}�,0�\>�1�z4G����k���={?��-��\����Z��w?����yԵ�,�wU�*��fC��]ᬓ,x[	K~:c䡬����s�� �2Q�k�3qpύe�=y�^uA� b�8S�(C��+�_ܶ}f��C�!��;�yo�|F��"Y��]/I�~���RN
ƻ� ���_u t�Sr�H*���&�_����T:�`Qg"�6���oG1w��VT6���{K���F�)�BĒ�s��gM�]<N�y��#���p�(%���Z�s'�G�t��<nRph���?��2c~�ۯ�ޠq$}}\��/>d�8}J����2}�U�H�("��s
��m� ���^jW�w���OF��DP�Q��a��cf7>9ۊ0̓uv�x��^��~�Hۢ:��'z��f[�f�5����dg��{���`TS�*9d������ݟ'�Lj��/����LlK'�����]"����ƢuZ�s��*;$�bo��jh�fw��qo��PD���z�j�t���c�;|H������,���2�a��Ж�C��kcĠ����z���a��#<Kq	O�J���7ZMR�|�t���g9a����y�XAҴ��̱�[�����y��|����lP�(]+���-�����Aʶ�<oC��z٭眤��8�������'Ց�lO@��׋�i�ÖB�^����BƼ5����}��{XU���m���jx��I�����6ȹU6�m���	�S>�J�����'�̨��zq]��r��J>#;��x��kk�[�o^�5��IQ��
�Ƚ���o��I�d'0h{>i����)��a��$!�k����@�����3 m���:/��*u��5��L�:���>ם���TD7\���(if�N��������J.MsZT�3e�P��	�K�8-��a�Xǲ.٥M����\�� �g��t�n��|�k�Ito�s*X�BQv��1����,A;.&>��"1a̱�%,��V�
�ю
�?�Q�,	T��N=���za�k�4_u�f�3��"�_9c��rp_0�([F�H��<l7X(^��ςg�ʹ���<~�H��9�xH� ����!y��d�&����+^���O'��G��� M��\�$Y��qɑ�9�϶ĀVS' �sUE[g�7�&brLQ̩g?���7�:)��gu����<���q�q��;hA��lE���T�-wg�|�}���������u���{��>���;x%dO�R�ց�g�6m�:{ќ?��m#��%r���G���SN�,���δ�<��R��k�� �N\^��S?���z��W�C�{V{�k����
�W����7�!ڭF���S:�Eq�|���s�SF�����d�,��<B*:��w�0��FI ��FJ5����_:Y�yl�3��ZX(��1�Pgՙ�ߗ{a+�<�[4��9�8|9�(E2R �����
Fk8��#�<����oɜ�bbd��r��F�Ń��F���j��v*��O�"��RZ]���1pC����
)礷fb�
D[�r�0�;.c����������"}_X$>6n͊�g܎������^��1ӄCY5�HI����q<T�� �_ݧ���X�"�=�;
�'��X�����<I
���ˡ����������2j\���(��9���eS�ytճZr��}z�"������MRΜ!O���m�(���a#��,Z
o�>��x�rMH�ÎòO[�f�ض^��_}�z56��o�pa��Nr�|n����R͸��
����F4�uO�ʘ`տ.xEc���Ra����-g���{�"���F�\e�+l]�۰�c*O1��b�[w�u�]2�۝�h��۶1xj8e]�\��V�V� �yBߩ�&L�s.�����%sd�C��fB��w�F@��I���x�u�}ŷɞr�c�7��qR�f���z���kjI3����oo�*�V�j����mB���v ��ڴ� s?������Be+�W���̄R�^Kq�����p�`��>e�xO�St���)P���׬�?I�<�^ ��)d��<%��@N�3��� ���[)���*�6j}�`-�ǲ�4��B�"�P���#�l�t��0k�_�_R��dM��_˲zf�M2��ٖ
c�@����ʑl�$����5�S@�k8�6��]}فR���n{@P���Jxۿ�Y:%j
V5��zryE���U|�4��@����b&y�AI���ھ�iM��Y,dۇ�+1����toI��ti����
�_]#y�ص<g���|[b���mF�����V3��c�ƪ���9�	��0ѓe�\�dJ�!��ݔﰩ��eo;���3�����ߠ�tA2��>����\�[�B�9K�m�(I�$�E�ru��4��4�K���"R�����ټ��f9�!����/�m�'�j�/�o�*�s<��y |�QM=�&���3u�J	��H����l�Lr��`2w1L�]"�7���Y4�'�u�֝�狹�Z��hM�p���y�~�c�b�{��>�ݶ,܆�`y6��"nP[��n��W�4d2��f9Oqy��:ؿ*�̃&�o�HT�𰴋*p���"��ps;����{��Zy��`�kEZ�,���?� C��1��m��c�n�5>A�� ��Ce�N>J����1�lg�����Y�jVeVYwP�p���r9/��Z<�7��g�o�9���n'���E1c*��ji�w�2�c����Ń�
��R�͉e
m���Ĥ�^Tg\4qaS�����MiQ{emѥ�x���0���%�7U�<J� ���DM>��SY��3ɀ�H9A�)!��;�v>��R�����&Ɛ�%��^���o|%��`���
�zw4c�R��h�*o�6�\����U�u"<2E�y�Xt��؞�Z�R37v��|�Q�4Ǽ
������|���qo�>�C�.^��ul�����J(��?�@�;�4�Ś�/p[8ۄ�����t
*�W).w6��b��������>�ohɏ7�!ʦt�t�j��G`�Z(z�pR����!�rj:k���=����� ^i���Ig����%�&��u�I۠�@�W{�o= zQYJ��E(��l���'�b^�?ʮ�~T�BH�����ED�t^��3��x≿�-]밺�9��q�'�#ܛ����+쐥>�'f l���?J�d����l�� %iۑ�&�����޷埩�/��o "5cfB�̍����]�
Rd��} �2����q?z0jT=�6a�?�6�߭�JT���}jr6w� [I ���4+��:r��{���dD>C�E���:u����Dg'�m��q-��!z���H��b�D�~��	�~�^�O�!fj��S0[A@��gMr=�F}�a����L&8NS��D���:ݻ�(��Y�f�$*��c�)m?i�@~�^�_\�Ċ����<��?µ�7/��x\ՠ���1����m2�'Ä{�n�L8:���dPhϰ�p[�[���]��RD��Z��Pr��äPl{���o�T<tl��T�'y^pՐ�6;{��=e,���Ƈ-r���RQ�27���1�X������A�	��+������_L�K��Ğdq.��mf�j�Ns�I���g�,=�%�R[�-�~��R��m+%��\G�J� bLn|��c[�!|D�}�tͮ�������Kf���C{�OG�m1��t�i��G&`|��i]k� �g�m����껙��5O�w�f�L�Er�ƬC0��X�j2ܖ)�e����lk�ۚ)8ы ��, �4B��)p��e�p�6�F�e�EH��=��P�3(QGIY]6�Q�S�xI5Ϛf���;�gׄҷ��h{z��� ҽ�Xc�zz��ɪ3( =�Y1ς�{e�V�eJ89u#�!�w�g�ӽѷ54F`�}�R�|������h�q�c��%�w|N�&85�U���W��q)�s|� uGM���Z��<�o0�f�X�A�?�e�b����)�x�6��\X�x�������x\3\��w,8V�_|�+�M,g��=�{V�q&k��#�.��i��т��$���M�j�c�:	�l����v�**�,>P�.7k�c��KT�1��w9E��`�!(���Qk$ۉVDt;Yp}%`��v�4�+���2vQ��4���7)��"��eqG���}�Z=��Z`��.(F�أ[�?ٱ�;ߊS&+�2�˰�Yoo���IQ��0<*6T� �q��y D�|���q<;�%"����g�����$~���Q���:���������D=2r�C�ЖO�蹱�W�$���IG=�\��ؗ��o�X)7������(>��i�/0i��x}t^��0E<tZ;,��@��#a�T�y{yB4��X��|0����;` �f?�M��J�>�⽹^&S��KH�D#\M���;�n3�}̷}m��t����x�#��M�=5��*}�ͦ��ɦ�� �as�@��8`��hwٚI�`��;{=�G#��]=�[�u����{5��+N;�a�[#��_@e^6f��T�����	�gna�!�Ab���o�f��#��A���̇��)��>�
�	�|��[{H�p`��ҢF5��[2Џ�Ȅ�i�U��mΗ�L�P�6������pT@�dZ���N�����4��,�����Y�M�p�+�B��8h�	]M�6��Y���tu5�:w�E���j6ĵ���[q���7����ڧ>\�$0��_e/ޭ��g��	rޱ��G�v�(��%�Ό��FE�&���H�Z�=�`�����}�yM�-�=�F��r:�`�H���Q�7����z9g�I��]��
�J���ǫz���L�)��S+Y�C{Ȕe�zY#�mS9t�[i�;2�c��{��V��E�̖5粷œ�p���φY�	�R���q�^���6�C��A�/�xо׏�~�?;/���kf&�Lc��`TZR�*67���ŋ:]&�����h�;�u�y��dȘe�EW�ɷ��K�kQ���brz��^K-!K&�����:�3��o78D𴹜�۬�dz6�y/N)�I�P��ߢ��҆{��Х�_ٖ�e�á�����/H��ϩ
	@����-e�T9�����"�Y��Gwv��w�J��b܏��{�����ە5�)�������!U�l�sDg	����ǲ�3��k���Ej723k3�U�ouR+��J��R�������~��y/�;#�q�i������#@u�G��KE��3]��`~����%G#dǴ���܂��e�&R��zR3���M��υ��aFj}����]AĶ-�k<zѓ���V��LXA:Y�^� �*��W�i�-����m'�5����Hk
~�=�Xp�6+bE9ṭg�t'C��&j����vc���s��K_4�8�mBU�,LEϕ0a?!jaM�b_�j�[��b�_��Թ9s���s�fYɤ�e��3�T�aL��������x�D	U�[�|�H�a�a����l=��i���.k|+�}������&x>|���5�Rr��h���B��}�Ss��eeB�O��CE�t�@yW��K9(%��z�	(i�|:������U���uɘ���b�7�w�;U�K�<|2"�aCT/-Sw�kE��� ,�IO���ϫn�4�Lɼ�?��lq'2XB�Oy�7��R��OgCa����Cf*�ݶE�$0���gL�E�چ��w蚍��=�L	3G��)���99���z���ӀG,�������sm�(�n�ۈK�S���H�����^��~c��ٝ�*�#|M}�)���=	Z�4����1�j��BO��P��;�VR�P�u�]�A�S����j��^El�q�.Խ�ۚ(|�t�K5$�}A����{�S���	%\����go@�#	���r?�9�ƈ�*�GX_��h�Q���jZ�|�W��M�׮ ��v�/R�v��u��N�����J�G�X�M�U�<i���ez��U;�vɪ��:�2pp��I���ᢘԭk��w���'�waao�F�j�@�����,���]��m-�M]	O�-�s�}��н�Pb�3@���=}͈-��iL�
]��z>�I!�Z"3�IR^NH�|�i�)S�vՅ��LC�����ZΈ��bʉ�Cl8���㸱�f�����1�?r�yF�c�pB5<\�#�ʯ��E3O�v���t�����rVf�����h�>B&�ƙ'I'�ӧߑE��4+m�)�MTV�2����>ݒzq�LC��C�P���`�Xh-����4�Oa��L��]��v	TEr�LbÖ��#)�X�Lp�㋾L�$6�ƴlx�����N�����9�;4�B��V�����h{�5�ډ�Pd���b�0�7�?S�1�\D��G�`ӂD �t%G�fS�u7(>=[-�zG���)Ⱦ|ޅ��l��a�E�<I�l�)���%XE��<���4p�Ik�M��V�p�d�OB��5y#G�>��.�Y��p�Aǁ���H�
d���w���M��fDH���:�g�$*`畄fYx���7STB��"�^���c��]�h��h�H'8@(���f��&%��B���u����W�Ir*����,ZSNҒ��-�}�z#2+uPeΊ�Q�#f�U����I�����ƃq�UH�C�<��yS�nQj����o�`��
�tSNI��2H��B�J}�����_9��7���I��F��q�6��!t�z 睫7��H��bI�~����-����-Y9��9}�[�8�}�ppK,<���N�m5G������\�k����8y+�fC���&��UE�~~�!R`�fw������StF� �;;����0��^R`��8�O�����v�y����*�.'9զ��� �S>rjF�󁴩�4��cC���������V<;а�;I�<� W��-C���"l�׳�%m�p�|�ݜv�Z���_�Ply���	OLN�Sav�~�7���ㇱ�������ĳ2�1��̉��P�B����-�S,���5E�
`/�S/�n�Z�S.��S�j�: ����'�OH� �FT��bS�[=����iba����~�8OD�c�p��)�єi�V3 ���<{�Ğ�-�Ia1�a��cG[�&���LH�|`]�nQ�������vܓ'l���$���v8�p�&�N4���� %��L��>S��I'C�����N�\}���U)Ĭ��7�n��g�*^A�6�9Nhd�Z!�E�ֆL5�`C�@��J\E�Jh2lN����y������be������'�T�Ŵ�~���B�5�vW��F3��f�"S-Սjp�v��N�"�f�X\�S������R�a�P�dJᤏO����~8D��B���	Q�d�
��N�ȳt�x�Ϗ'ː8���� ��3�h�UYo�zT��m{>�tR�ڹ�C�m,Rc
?[���2
�u���&���.OG�����N`�p~�U���$ǆN�s;8M�v<��G�{�0�\&Hn�cR�NuZ&��9�3���`�1]DS���s/el�����+y!D{�2W�S��S�����1"�-����Z��.�q�����3�LSBÀ@Gb��><��[W�i3������SKZZ��� �	vM��N���Á��]�߶�Z�H����N��>�js��=4˱��|d���mS��|��U��8<�[�jB��4� �!��uȣ��>�K��k���8����l��J#w��'ݿ�Q[_�(�/4�1a�4)<Ϡ�F�C�-,+�}�`KV&Kc�̧8W���u���z;^�5<N�z�7�K��a_;�u��e���y����k��\��������]��&z<}Z�*k����\��b�?kMF����R�C�6��I,�gګ��ɡ%�>��~�@R%�n&m�l0Q ��q���͠�
Т���O���͘���G�K�B˰zƗy�~�>R�by!�I3LC���Ƚ�9|4AL��=ėқ(��Uބ��05�X(�ȉ1��.n��M�)�����J�%�4�+TCF�B�/�~ R➺�fa/�Ki�X��-���D�ߗua�
9��	TyF��_f	���@/y+3^��=�Bt����7Ї�q�j�)�����0�J�����X�F\=iQnd�HWjGr-T��ne
V��á�a6`��q|r<b>3D�����n{������j��D���i��go\?z���]���p��8���a�۾��`[o���|9QZ!��۔����;��5�]�פ"��C�k�����a�8Qބ��\��uw�\Ev���5#�N:�l�M���}��0�%.?ñN�(�u�T�.� Y�t���"��\����։�-�`�����^���z��m�"�w܌�xq�E�_��a���̯�}�&��-�N���0Eqq�L-�``M�:�7�^��J�k�����z��b%k��`Wo!3@�,�0��f�P%�\n�V��V���ue�~;���)b'�tZ1V�Wn1��=�.3����:1!��ݨmn��<��(T�����6d��In'��?�υ���$J�����8��"�V�0��`�'��B�N(-8T�i�{���=Z�쎮�4>Y�(dPh��Jڦ#E�ŀB���o�r[�\np{�^���b��Q�=g�B`��ŷ<m�@���	�����P�	2�_�i�	q���9��/�a���_�O�|1�H�{d 㩺�5&�����Z�����sP��r�n�umYPkk]�+��<>䁟{�����ty���2����uV0��#�R��Vu�����ݮ�ڿF�WE�dVbv��]|}�'�=!$�������n��}W����:�{ijz&�� ]�)jv�2��&rMOb��Y��;�]���%��P�2�:&D����G3�,F���G�;p�r;�w��ga7�����U��ˇ�^[T���S��S1� �8��)M�� gU��V�p���A��,.��d���)h�v*A�Ѽ|w6c'2��,g��%�9)M�Z?�ּoi��6�%�W9������^ګd~r��D���X�������9�Ͱ���~}��n#���AG*S���(�.��,��#������E�H�aS�3x2�J'�-���q7��æ��pi;�� �@A����O�S���ON�<�u�-��]rX+c���8)��Iٻ@����l�
�1��s�=682EԓHX)h�����a�;��wW�K9U�2��-���T[z��ec����8�7�8���#(�G�*���qB ��R*���#!��P(
u��S�dǽ̸5��~�o}<Z��I����I�jJ=��"�T�zĢAK�g�;xG%�͓ּ��{w�I��b{'x:/W#>�å�t�a��s���˦��]U��y֎�A�A�`�-�)��[:	��!>�m뉒 �=I��*�Ș$���e�f�Zהڐ�]z��T0�t���#xy�7���c�^q��؎�sW*L�g���vU]v%��ш��hU���1�8ֿV;M�S,����!?q�C�F��B���W{�^T> ���on��Qe�M:�����h�c\��/</Ic2$���[�Y��P�#�a�DtR�Ѓ�����M`�-4��$���~�MvH������q	oD���M㞥�
�M��283�Cd�� ��RZ��#����a�]ˈe?�l��#�<ś�-��.����J�Zq�N���{Y����#pD�10�����)m�dt.���w����`2Ldn�
����X�u�ut���`,Z��/^z��=k��B'	���W{y/��A[',�Yx��/�q���Ә6R �nt�p���ѹ	Xr�ۅ`^�&a�`�7*���wGǕ$�FSݮ���>��2۬�c#�-0���;��3��S��-S�LX	G���-�5)�s�3�fiU.w��'�p�]F��3�H���c�>�O�#LK0��ޟ��.,�ֿS�^��h�?�wD�9�pTe��z���8)V�����i����l�g ����`�̭a!>��~^�WY6i�ِۨ(����[)�.��n��LTqsAj��Xo?��Q�(���>S����l'��{hX��+�8:o�8������	��8~��l���^���~v�j�w��2A�� O��sM���޷�~����|8Z�A�r#�'x�����tg�-&�(B���^�т�d�Z&T����4�몎"�p,\�M��LSZ3JUU�sh���4x �k�F��XQ�~pL_1��0s7|HR��� ��X�A>�l���q%7W���2��oʺV�D��]����d���ٔY<���gg�5oМ�L@2�`vP=�/��V-U0��:�iE+��Ċe�K�����|#v���A1�����BKY+:p��&C$��3aw��o^��w�j���:`�±���>+<oC:k0AjS�V#�	�i����S��\���J��"l������`���U�|K�� ,ʂ3"��������3sw�s	�
4{�Bs�A�T���0�n{d.p��dA!}=gz`%(�P?1��!�ł�C'�i|�0p快��j�%X���}�h*sBO�8��؁�6�����I$t)W��I*��qP�ڿџ`4�ڷ�;R��1�t�j8ߕ����4aJ#��NC	I���	�~���������ZRk;�DEk�F��ȩ�T4;�m/�����a3��a?A�}w  fc�����KOPa��Jĝ��I�?:3G+9���"דnNM�L"{���ڒv.Up���FqŊT�)?Q�HTx�F �;���q����� 9�p%-��1 ��2��Q�1�!���2��V\�h�E�`#��#0�е~�����G���:��>����o��k0��� eV1'����T�������O(n�߽��7XE�7[��I#�'�Rx&0]��L�O�������BU�z.4�q�/���B\=\��}TGa�]5���iѽP�?qn�+��b�IU��KU,� �)�Ftw�U�T�:�W"ߐ:��b�..+�Z+A�E��>���d>�u��.�\�c�
��ܪ�Wt�)�#rh�T��vbr�B ��ə�y�0q���`@M�"�b�g@;a���/�h�]�k���	��7D��Ľ�ĥ�6�4�W��=��T�WS�j����4��_�G<%�A>!s��W��%2E����.E�f���Ձ�CTG����q	�_I��� �b M�8.��h��tZGV[e4][H���l~)
.+��$�.�K+�1�xs���^���ދ�!y�}_��=�6i�J��y��կ_g�zF�Z��p��h_ �sJ�6��P��K4�3/ɱ�ڰQ*9e��K�hm ��i� 9m�H@^|��\tR�k�	��"]3�㆟;)�J�o˥�Ҟ����[�9�oɹ��q�1����K����I��1�`ͩX�(�=��v_�0
��/*�p!̨ދ�.���Սg��2#�qDԿ�.�S�G M/7Ov��~c��о��q"=��]=>�bK_�ɯD J];�ʭHic���J�kbz�O>d��u�!'u܂�}�F{w��y���!�{U����O�~Е���g�gW]&��gc(�Ñ�+�Aڈͳ'��*��M�X `��	�E�I�٤�OI�J��j�&�lņ����,���f��a����J�)s�wN�˿����o�f���}���8l)��*V(�0�K�oا,c-u1��ɾ�E r��غʎ�K��@'\�Q�C}U��b�n;�W�]���dD�t�=u��D�3��5�����;��/�ռ�K�V�O�%B\��H��;��硆�J�s<j[ZuV'�6$����}5n\�y�_���s��uhgN_m~�L3>Za�I���6��R4;���m4�}�� �tBd4h�)aqg�3Z6�P"0������R�=�ěX�+�=�	���LO�θ�e�`A2�u���/]HE�8������lY���/XN;�r9�T\3wWG+.��G�"��#4��&��I�߫�������4�hO�,���T47;�u&S��!�]��݀�х(	�G�vT��������Mj$k��O�"d�r���N9�����W�JA �^��j��ؔ�)I�1$r`G�5��@ <��l�R"��E�p~�[_�G�O�k[���e,�k!A�i+BL\�������!�_�Oa�S���ZQi�U�s� {;A<���U'C�Vpt��i"�e�Oe1�����FF��}��.ap�z���L���g�L�Z�\Dʺ�j����������!ئ�ڈ$�ֵja���\���tT� �a����47�@;�=@�K�~lm��%���IѬ�����f� �/���<%H��7ؼ�M$�˗�/��+ ?D�BKB��x}FJ�{���etVN�m��n�mا�v��8�CS����X�h�|�MF8o ��N'�sq�!'Ѳ��b�	����(�lK�11�9��D���B��:c͑ye�5ؽ��{�"4���2�@�
6w�/"�o��w4��Ƣ E̦���(�G�z�m�C�P��<!��J춦���=(���
�Ȣ˩�w��jf6pF؟G`�dR��`��T���q<ߙ�J����)rιd�Ǯ8�c����5Z���{�c���" �V�T��ں�r��{h r^`��S�w��z���L�5��'l^��ᗡ�<$�@~��|.���)�>������#��i�:�f�vƙ�ӗ=�l��&>d78W���G�=��;'��AT�X�5����((�Y^;��[�<_]r�Th"N}�F.���]ym�Y�y�0�9K��,��z��N!����5�л�}��v���F���g�{�%���������!�J�����H\��H&!�Z��f�í����ߊ}�p���"���RU�3!��ǜJ�F�yIK��4�0��pG�c{Oy�)�L6���h���l���7w� ���g���ұ�I�~����*B}I�5��s2d�vh�#��Oܼ��y��ř��v�G��h��^E�B����t�-$�Y/̱Q��S�%��O�/��j��|k��튺�[W5��D��jvЅ�"3b��[�Rv��d֍[ �C8l{h�+?/	O�&�J��B�FӲ�s�+1������FȢ ���3�Z<>�PޠNl�Cr�e_��6o����S�+D'�X��J��?'B���9'b�}mxR����l����B�߆eh���D"�J���\�8`�f�V����!�m�L\�m�d�y>B�?�5i��U��bv;�5K<R�7࿹t���6���%�1�oT�j���<���WHz&1X�1T&�b�+{���5B
�=&e
�$�l+�//h�-fn�0�?��Q�N�t����ճv|���!�Y�k� ��Zhh�s�s6[�t�������X^ſ}�o��q~Z-��/5]
������b�yx(��� ��O��$��z8ٱ<��%�`.�)�eǧ�q����
v���϶�|�A&�� &��6�~ѳL��V�%���d�WB1�D���8f���Ugo�/��'�%�1U�=�7q��ݙO�0�|��l����Ѿ�.�sCMXNNdL����bje�V���yܡӇ�DbqLnh~`�&�L� �$��mn�q>��/�T ^r�C.�M�`w��z6�>����=�oQ�KSU�c��n�*ƍI��&#+�/)<�7`Tgg�*�D��wLV���J��$��K�l�����(<6�jlV�C]�����[�ʚ���QKފ`����'�hў�Q�$�cv������Wi7����<�J��f�2�'ca�������LM�N�/V�S���3k�E\K�ٱ5�oBF�X�ɛL��@��%`���(�ߑM7.@H��L/��	�v�x�R����>����)L�j��r}&�<�b���F�����<t�AN~^�(w+� &|�1���Ê�����-Z;�ߋ��3�0�HS��'�Y��`�DD�� r�ɕ,d�d��写�΀��n�*9���L̘v!���A�
��l���!3;Μ�j��-�}��R��)�'�=����gx�;�.> �I��R��6�Ë����Ց�U�����S�9]��qp0� wm�aQ�ٞ�݅d7"�ݾ��|��Z��� @w�>�%��tl�@��ȋ�HU�Z�zv�GC;��[��U�vԃ���q)d�m6���Ez_�&�v�7��X��l
��.O�3���юV��&x�]����)�<Js��z���N$�9����I��8a�V�/���s�8���(Y�c��P-�i�"�V����*�|S�Z*��RJY�Uɬ=&V��6.�����6.����.���h{����%H�$v@/KF�U�j�����a���H$?�M�e�:}%�T*��� �@��pgjc� <ؾr��G�A8eq\�>+�RN��[�[�a]��Ҵ<���-&�Iw����f����'9Ϻ�Wm�i��šׇ����G_�o	#�Ϩ1IF��~t@��2x�	�}Ҁ���	�B�S�$��ރ��3*k!�v�h��?y�c��R���=����3+I�B�X1�����Ym����;7�2�J�E.&��g���{Ҧ�:���BN	o�"�yE�O��7�'G0x���G79M�Z��F�s�望���0# 73���߆+ذM��/}���%Fo�1���o��% �*T�֪k��1� ��2aJ��s7҆�0xq�Q0�#��4�L�[>�>N&�﫠�Ǩ�A����">��з�c�;�eb
+6{��to�5������s�&ZRx���F��w��/�!�+�@P��3>�>g�6:�X�G?��HY󒑘E)�8����k�<y�PF%J	�<%�~��9�[1�H�<�Q`�Ux���I�
x��X���Q���na4#�C�e���B�W!��0��K6\�����m���s'�p.�Y_34?��'���*r�G�+�]4���u��k����p���h89t����@�(��!*|��"dL|?�>���6 ��t�a���	����G���!X�
s'� n�~1e�	�ҩAx��oݽf31�!,<�8ԶN��i��Ŧ]���k}���� �_a�3��f�	U��B&��C�鏽*C��8�a[ y)�g��ƑDǏ{�HѕXC��K����]�CS�Nziɥo$=N�O"�B�ut�#���7�N%5Ofm#�Wa�.j�ෟ��Á-��Hĳ���Q��������Ao�3jbY�T�s���c��o;�p����I����%��h�3g���R@����9m� :�0�@("����� ��"�|�<MFC\��2�{���)�o}�Ԇg���� � R���p�<�[���K7 f�+]�6g��/�v�`����>W\B���x~W	6���.�$0�0�6��>����&$spI��f$z��y�ZHz��u3K��P��oR=N4��p��.P�]�cZ$ix\���]د8��ZK�q8�淂�$.���� [,%f��bh����͕zz;��e������At3�hrܫ9qr�2R�om���͈�����6j���<�����6��֋}ڙ�/pJ�{�K��ݧ*u���΄�CL���MH@���H\���M�m����3�sOi�
�iX�?v#�~�V��<��鰠�����QCQc<���9��5Du.G͸'��w���(��q_َ��L
��de���]����j)(P��GA$�p"� ndF7�q�yl�0f��΋��V�R�񓱀�vo�vm��	u�1T�ƀ��y\.�~+4���#r��R� Piuۨ�Fe
Im�.x�)Xko���x���2�U\�`4�������A���O���΄��-�%��M����)�R�X((C�����\(�������H�[�[鶬g�
?��{��n����e!����%9��{��iͤBi
�[U�}��b�ȹ��`:"N�čL���&�8 ���Կ+k�{D_�gƢN���J�)��ȝ�����:��K�u|i)��2&�A^���L�6&�1�j��<5�욚�������+Ѵ��	5w�%K^�AN�"���H:�^~�e��(U�!�˗;N>���dh���rz�=E���N<���)U~*��"�[Ct��m [�J�KY�4�l�{\�bR��Ƥ���t��t���xH>���]lq�n1��'/݄��A�Dqx�2��Mö(	��R?���5���2��Ƹ��l��j��i�K���8��+@�..�ya]$�1��L{�K���_�G �2��4���!�1i%���E.�A�"���
�L��q]Juy&�.�h��s|.�v=,�,��бAD�W�6�[4�N]�L�#)=F�m]�5;;P�SF�Β���O`�3�H;p��y��^Ȍ�>��V�7�B���+���Z�Ƽ:����e^�8;�[�>$��;�fK|�U����hag�Rܙ[ڐ��\���S�53<4 �bB�?{0��64��<Ar��B6ƞ�
]]Xa#(OU�����T)z��I��&[�G��gpv</���$�43����t-���s��<܌1�	Imy�8����r'̯(k���Bg�t��x�Z��\+�tA�)������+�IID�~0�Wz�k�|l'9�`J�Oe��c��w�'�d�d���j	��msYACsʺ�+2�7 GLP���W<ש �9F�-� ��R��
�Vd�4v���z��_>'��a��V9tt��n�+|'r�������X\	ݨ�G��>�u�gd������ ��Hpl�{�*�+��`�y T�GP]��:O��F��!	��U��kר��o~�U��vyu}���M�kD��؈u���g�d�8�v��w�.��������^�u6(���ar#���me��3pt)�?x= ׿��5-�`v�o�7�%ݸ���S�6�eha���qt����WS	tBx��S�/,(������L`*y9s[j�TR���b�kTs@;&��J���4�NٔOJ���F|�	�ܵ��o���M,�Z��uP���	��\�#2kW��T�Q\e2��J�+��H��@O�(��`�eբ��(���^��&� ��IoD�(���#��|b!Y��y�J��ѕL�\���ޮ1`,���Ɖ�q���Ŀ̾h^����1^�-�]=�����!�)�C���1�
I^J�b��9:���6χ#������ ��"Y�M`�iӍ,*��:�|��4�n�._(�gT���N{NXO,�Mo�����@'.����'�����r��k��M��։��vި�w=~X����@;v�� ]��S�c�o���@�v��q���6'k,rZP�m�_��yb�{���B�2Ϝ���NC�T�9/�n�o�O`���F�-C�+j؝V�ݍ�О�'���ɻ M�mx��!
�ӆ2o}S�'R�}�E;���ħ���uh/eC�9*�������	����)��(3���?�'�����"��;!�`	�
�K���0�-��Dg��̌�3HH���*W0�윛���*54�|#x.��<H��]�u���c��l��A��!���xc�R
D	X+r�*@{�v��7���B�M�@��\��4����~ox������:6�:Ñ����
X��Pw�����?H����6&O�J����q�j*@��f�WXt�fI�t'@��'��r��J]�w�v�T�Zn���Z��b��pK�K�Љ����;����O�I�?�r1'�r}�&E�@2�*�!�8��=W�
$�����R�c�u!Ь��$�܄ۼ�Bb�g�N�j�F��x���}�ZvHU��a�36�m��Of�.n#pʴ�"�K���Z]Äh%�ڳ�^�cs�	aR/�k�T�}�f�]>���L��7گ�,��JŜ����?{~?��EzH&$�o����)���LMoT����@°���G�p�?2!S�M�d�Ya��4f�[J1ɦ�7��=l���S�Ŋ4�2�|�J�+U�;Iك/7͋j,�9 ���JP���%W�q����jD��Nv�)0*:\�#�]�hs8�8T��&�0RqRC�{�nX��C|fo�s;�-b\�2��q�&�ţ����H.�U�������K�I�,�9]m��2]jG�k�o���[��Jv�% ��R"���"��RtE���X�+s�u�(̞���z��Уq�� �l�q�l�ު��$�w�9QՋ$l�3X�C�5�GQ)��e�=DX��z1*��X_n���0����
�1_1������VY�5<A �W��q������E����*��"��oOx����/�MS{Ӱ	��f7���KP��u���+�
&Qw�E� zX��>	���Ɵ�t��������ȱY�霠���:�Z�~�����3��q���v.9��m�<�!��,vҠIm]8���A��z�`�}�a��8~�LɄ:��i;hNY;8�:O���|��$V6�|��+��;?�V�i���T edi|��'S�5��H�8�ŪƝ�{k�J���Y�f��-�k}����Y�S��Q��'(F�v�<��jd*�����2<��ZH��z��9����j��~�]��at}����$:�^A�s���6�*p{u�_S����ͣ;㟂�����eb�'<`�����ls��<�o���A��������[� ��d�֜Y�+�gI�l����	��'�QZg^yG/t����If�� ��F&��\IM[	4/�:��J��NTqe	������)ILP@�� !ɝ�Ɓ�u��A��N��j7W�zyh{�}C����0�:bls�����t~��5<c�DVN^�R���@ ��'K=@�5ַIk-;B���'��S^8�G$3� \*Z����c\��l���ڌ J��-��n��
���ո��y�7>�k������.b6x���!(}�A�f�7ǀ�p&�E���Di��h��?��"�Q~�^;W,��H6�@q21� ��[+�1XЫ^K�yMc?d̩�j}��|Rh�k�閯�5K�w�T��2I�ƅ�$��[B"Tc�Լ��{�BZ�'x��H3y�g�
��`͘��_}XbI[��߷uwP�E<����~gf\J�A�"�)L�d�iP���Ki�������P��^��S�H���|�6sb
ӻCF�@�I��ҥC����|(z��?�H�~���4�^���v9����𚗿╅�xYn2���V�N$�m���?K[����,���,�tVnO"����[���D�#f�BW��Z�޸�rj����:.N;W�b�G� K�+_?��5�o�=���:��#o������e\B�*B`6�n Tdb�3S^�|���d:�_�6��M�8\��]7�����i��9s��2�X�B�{u�֑֩�~�|D�'��������cdKn�J��h\�3���ܡ�����@$�
��G�)m�RVl�عh̖L�dm�Q�i��+��'����B���ҩ؄a	�˶�I�>@ǜeZ^+>�u��NX�;3Q��js��
c����i5�e2��F����m�$xWvdV�t�.5�k�ݓ%+�;P��c6��.���_K��iOc�H̙�6���㋗�*�~16�N��}������:�ܒ�(0��z��<vOP󧍠BH���4��%��k��g�LO+/�CZ�cL�>�d��5���N�(A��L7~�6qī�"��*y�޳7����M�(�<��]]�v�#����ٜ��[�a�&n��a�gV�9WE��VO^۵�W��/�]�K�S�Bo�߻$(�e^�L��H'����x��R�'�u���hR��@�p�nj0�*=��� QR��Ԡ��,�-/>w�Ėq]�=E!���ƹ�.9��[l�̴�I�cWށA3��"�/=O�v��(�o��p���y���Ԙփ�.@W�`�B-	ي����8y����ro�����'Cv�3�B�J)��(�mw�]�~|�dl���2+��M E1Y�a��n�"�їk���Y��@�Q;6o�to����;hO���p��{�w�O;��:&֘�;q�_nuظCi��ig���H�2Xe>ݒ��y�ܟ1�(�AE�1�����)z wq�ҭo��y��=�Eh���㐫�vx�c۳�U�MlEX�h`��׆M�aq3T��S �G�\���0w�s�W�Z�ٙR{�-])�,�o��#s,�Mw��N�l��x�q~ś�]� �oP���Qσ�[�����e�s���VQ�4-*�=2z�[/:�1T���i�/��"�}��R�2�^�,��8����'��!g��8=(x*<��_Y��l��AQ�ar��yT-��\�i��שm �.�P��׊[�N�!�3O�eZM�C�O��kS�9��*S�7�d-:��>s>g?TfJ��c�ILЛ2��H{������H�v�!.&2 J�Y )�
�_ޮ@.�M��;ٽHr`W5�-�X��޼G����ae�����p��=���m"ȗ���b{z�Ø	S0SF��b럢
R°�84�p�3�%����g�O�S�Y�9�u��%2�(��R����G�ٸ@x�r�~�Qi+F���X:ɝ�侃�c�{�ޓt��9O�.E�# Y��R�}��`�i^ݐ�f�3p�c�-�1Uv�����5�\M��bʶ��6d bI�2�І'�EѬ�;��5+��>i��R���F�}q��&��"t�&�;��:`���?ߪr�z�A_�����5zH��9��BE�i�f[P�F߭�����H�|={1K����6�.�"فs1�2��;"Z�'�q���aye��wPu͚Хm�T���54x�
�$�J޼(zBa�������'-�.F'�!���al�c�{�{�}A�q�F�C�U#
m�(��$�QRZ�B	JRFJfA�ዉciS-�%�bX˷��E��,8���t�4CL:kO�D�N��2?�'_l˚G��)qw��+&��eg��ƌ]Su��)�bL<�����B��t�39$4	ok�	A:���2�=������O�CN�V*�l�@wޞ��>����ٙ\=�J{9S�{�!Uo�8N�x̹���m��i�y+�c㡮����a���x5Y��Uc�I��]�g7�>:c�KM��%�(\���浓��o���s�2<��LEx�0oɓ�v�)o��6�ܟ|e-�����5�T�B���ƃF�Y��}>���KY�u����<�=Of�M�^��s��C���+sb����om���!~�6���p4T�_ʙ��w����o�V��ݜR|�~��&���f�AOf����0��nL���@�_��Z ��̬"8S��L;�⾒�ו5��������(���y�O+ڕ�F�/���gN�H|RA,oF��
����Y��IC
X��D�=x�cv�����n53q��X{���D��"�x���R\���jg#�h��Ul�G��P�,e�u{�I�ʓ���*z�������Χ�z���6�����-F�Y�k�}n�h��y� 6�j�ظ=.i��SJ�Y���e�yB�m�L�oɗ�+�}U�bl��sN�6m�r�H5I���ʳY��b�_e����1ܯ�}���{���O�����*U'�w���$�5DM��	Xvt�NW
���o��P����~T�@%�mM6�ޅ�8�͍4vlBr�=	���>�9$H��G�HD�\���`�U%4@� ���|rwߘ�{m�i&�O������AT����p@�77.�V�P���Z,q��b/��X�g�6@5v��z�E���' i�<X��t ��ל���4,��I&�g�P�0�zd��i@�Er|�F5�duf�M�y_������.D�p�����ɜh�j�0��������!Hn��x��L���X���L��
 Q�U�u��S�|es��8�#��&S3�
)�Wcޮ���C9�ޭ�F�dwx��%�8@l�BR1Ӌ�	����/;��3��:�p�ьz�]�N�>Ш�|5�e���j�-#|��,uXUt={+��y(�;/٬I�(��F�[Sh�o�kd,��L�ؠ�T�}Y��3Y}�G� �F��H������"��� 9�m�����Y�%��MA� ��m�;3�dӿ�/���W���uWK�Zh�i d��d�	1�BO\�Q�n�!�C�'������M
���]�NQ�C��fhZL-Z!m��$�כY=ng���\��*���ʷ]{�Ĵ�����F�"��� �n#����l� h�&��TD˥V��U�9��}�����(X�)��<�P)Ŵ?���߻k��x�ܽ�|���,��$�	<��k�ן�}��(@�D�%O����y;.�QD?�0⨂_��wJ"�F�{�E���R���!�|La�<ei�&�}Hp��r?���tJ�8���v2:`*��쵈9���R�v����0��L��g&d�V~|� ?!"M��G�zڱ�
%��gu��г��:�Pئ�%tQ���V�CU�y#F�3��̩�/��j�B��?A�Z<e+y��*�O��k&���i�n�C:Ō��zg�6�ݥ��,�'Al.�����\�+���G?�7��њ���o�ke�%^����֚�˶o?NZ���/lͪ�dRu�RyY��N��S/�ʵN:�U��JiLۏS�ͧ}$�Z��2>/F���w >|��ܿlY�m}ǜ׏r	�)��E��Ϥ�=~�cElÁ���dVq��ڳ*d�d.=�?z�L?`����,�ϫE�H�ᎁ��F�I$�� �c^T�̓Gcu��	����!Al�a��FTڐ���׏�/��<�_2�[-�w�U*��*\P�Nޔ��`���\�~B�Y�K��GT@�ǻJY��DQ2U)�'�H9?qYg�t������㼄��+�$cO��oH� ~�m�mãw��)&b*Y�� 6`L��OP�qpl�RDu��C���iD�05���-��}\��*�z:I�h�f�����J��h]*�����@��𩴙���+�qύ��J�ғJϯ�B�ɔ1���$���%��i�a`Q�X���3d7T/�B���a�˛@0�X<Ǎv�L�&p|]i3kA�i?���?0vP�G��lS�����jZ��5�{��ܵ}�-~ә<�FR��B�һZj�XO����aI�߄�'��@�Qr浝�R���ɡ*=q$��j�VIb\Uۃ��=�|�`�x��?��:L���Ұ�2�#�͸(���y���΅�0����ʷ�U�b��Z�=�5�.��[�ë+	f_G�ض��6Ud9X$������:?Â�-�Hߴ��WR�0�.m��%ۏ��O-�~�ӝ���Z�2�wӟ��PO��t�R
�5��$�p`}��(� &cd�o��sqIO�w��!}�=jɃ9��i�=����M�w�����4�_^�$��t�e�Mk�ו�e{`ZܓC+�2��2.}h	�޾zߘ�(�?��6��He���ħ����jq��E��4)G���ʳt�M��-/�ZCV*mߖ�ږ���R�F����,�:�qe�໵s����7xhe�8� ��V60�(���t(�F�Y8��h�e�<,{��,ݬ1Gbʚ��uy�1#UW֧�\�����R��Զ�����Co���쾸G�h���j�+%���2?��?$��{�raR�.AJ�t)�g������g��i��O�YKE��̏��Jq���c�noA9��I�^�U"Y�!�ri�U�B�1͞�����}�H�t0���!�ڄ�ԙ�M4n*�H�d"2�F��k�Bj�E=8ῷ���f��>sO+1�v�e�,lek9C�B� ܩ�w��}t�;)E�8)�<�M2$Y��=�Зߢ�aX��3*"�����HHs��!%z�B��G���0�m��*|��O)y��*�`�L�#-�0�]o���E3�?Jݽ�r�
�^ɸ���T�8���V��>�qd?�U�ygWz�0��G�~��� ���@�s�e�Wsd̳b*��
��Ͱ�*���Gښ��/6��Jٶ,8`�xqY�0��5�TT\֚��43��K� ����I<EZ4���j8��^_�웝�h*��D��:$~Lx.�����J����&�/)-˰��.E�}�-C�)��W��`jU#/�S�h����o���?*2��!��s[}�LЂ8�_9$�cXxakh�������e���3����R��S��w\�2)%4ځ nynX�6�+<��nme���S���$���EE� �r:���dm�b��r���e�P��Y)�Pl��bHkx���$�ּ6?>��^�v�.�D=b�ֱMcÄͼ�*OD<�h���;%pZ�#�i�B��Nr�D�0Ъ?���ťQ�l��'QHt��u����1ނu<��$�έ݉TZNӍc L�و��[�nIy�0��l{���ö�������xG�Ӧ�����zM��q#`Ι!�%wK��لTa����q}*�q������C�;�G�C� �j���
�`��m�������2�q`W�0���-xRiހ5k'��	�NN&�#6������ˣç�t��񲤩�B��� �v_�j��j �0a>���V�n8�Gd��ʊݢ� ��<uF�ns��*7�*�Dz��A��t���¬D&x�.���-�~��ݐ%�1�_�p��
C!:�;��{���4C�I��{�w���o�}�Q�����K��R�O�k�,O��������7�#�F̸���w!��I���f���^1-�*B��)�<(�����]
����%-���OI���d�H�񀢮`=�h�z�n-gK��)^A%�jJ��Pw�q�������c6�T�T���*r���|�P����B�݈/ �Dp�v��1�Ui&Y�j�6#|w�6��dC7��S�#[�kI,�����[+���>v�*��$;1cۑ�Q��pvA�F���; L"I��ȶ��1�ͪ�ˡ{l���i�ߩA�28:q�7���G����w6�s�6f:�zP�),zDq�%�Wb�%�Vǖ��Z��[��/��^�b�G���5�V�t_��=;�9�5��B�@����a�w�m��ٻ� �Zr�H0�������/fش�J��h[�6�*�jp�hi���)���	�M�=��q���g��c���04<cw('O�"��wC�̊�mkZP2�`�O���	`�0����Q_ȇvP)��F�vk�@�Do
t��!&��('ϸ�c��9�����5%����>_���=�aM�"�S�5E���J"���ұ��A�y���������"����w�� &QY"^�3�GV��?��'�L
\�����	~��7|o�c
8�E�p�h�����d|�5��i��Z��6�U�&O@����a��'n�(�P��h^PA�!����t@�]M�Zt��Fe<X�x�C��l�J��,0	2$�|�	N�	�S����p�E�������[��4���휳q$g���AD���h}G�sFը-�<��+���?N��ӎ�I�j��P�l2����d/K�3�-�%�\��ȵ ��˧�y	W�Aa��y���N=7���`Sh�ll�n�"wk��RJ&�vP���W�h�by��C�tԅԱ��ES�К
[l��1��_���]a��T�8F ���<�!_1資g���b�wtU{��	�l�N~4�Y�qMȸ���+��*7j�+�a�DtrjTwy���`r�4_�d�WF@�'4�A�+��}��,�zB��������Q~�W��qU2�g��Ӽʙ��+=+�X鯒A����l֏�Mx��ꦑ����(cޠע�GBVɎ���M��y׎S)��Y��Xb��PU�q�$l��<R=�b˯�G���I4� 𬟴"'h9�E�������=A��[i�\��x���`6�O�O��͈6{eJfH1"�x4���L�+c�<J�)2�x�4f^�/j�Qn���J�<"~�>��l�֔�K�]��-��*/�F��5���@�<if%�L^7E+ِ�t'C�r��P�z���Uz�[W����c�t"2m1�$���ˇ=��Q�:�5��pkB�.]}���Q	����H����Spsf���|��el�&/g��7��*JX� @#���w���H�1�^�(l)n�MsO����sN������u\8;��>����lP�~	?$	��9K�4�/6գVa�;ǋ�w�t8���a0M�i�@E���څe��|�0�s��4[w\�)�^�쑵IqC�6�sUe&.���g����6R����E�|��\%')i<����v��(��}�I��n_v�u�٨����QwT�m�Ps
����Vh�H�仡�=:v��Ph���RӦE���3Jb�\�&�,Ѻ37��gğ�eY�3��1��~�&���3�dH\Q�hn��G��i��F��9e��y�.��jo&�-=�Iy(G��Q?�4ee����_����%V�D�g��(����e�f�nu��P���9FL%ʂ�m����*���h떄MQ���nCk�Xq~��⟈��D�@�V���-f"ٱ��$�}���4$�Z&�j�L�$�>�&edH=��~F=|kX	��lQ�z��]˶kPbA"76᠃P�к��g���6