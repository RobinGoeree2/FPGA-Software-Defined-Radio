��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏����⽸���D��6T�8�{N�/i�kf�!�6��̋"X��:�����\N(h�-����}!���1�����4�0���S��k��Xd�d���{�8�%���AHǚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|/K�^!�� �Ϊ�I.F3�h�]D���� �1x�ϓ�k�K]b�ec���9�̑�2�۰�}EW��E�aǧ�b��S��+�/Aė �d��׫�~^^��y�4�4pjTK��~<OS[�EI|�ݾ�wi���tW3|��.�O���u�E`��C�g�"�~��~�<�@{�<��Nּ��~�K5��o�=�^*����q_�u�~�#��*��Yd��77�U9t) ):i��6�"���B"�3��`��4E�pI �jpRxDB�-}/9I�Fn���K�TW?�7J�����~��Mg�QʭO�E�x l���T���-�/K8֑2E?�����*�ݞ�1�4-!��U��=/���,C|ͼ׆���.��K�N�=��F�;m�\����T�[���?��=i�}Y_3�%]k��'�HA���g�$�4�j�}����Q׳��}E'b��g�}�;�CW�6
�����f�H���4�_!= �	����)`����A��Z*S^�������R��eXx�z�L�$�q��ɫ}�ڷa�;�θψ�t��՗Z���=/P�v]D�����+(xۀ���^ �e��1E�&ȓx�DE����U�/��]I�V2i���f��A<�>�}t�XJ�$`7���ٜ��9AЌ���'�n�k�M��D�� �P�9����6�%{Y��|鯲��Rt������l(E�G1�l�{A��J���͆q�k���\wɋ�G�<�b.�8������j�C�-TF>����H`���M�g�OR@- k�k���r_�<���sPy>[/����F�Me���\��������G"�v�F#�ę4���RUz�MGz���`�����t��
"�O��	�{D�|@h�dة<b��҆zF�_�6������7�������l����`͸#�^/ȡ�u�	|'<#S(�C��/�*S�K�&�9�yO���R����d
�����n��lv��L�l��A\�؀H�>� '�i_�5�T�@Fʩ�¹̄6��S�c	�\�Β�!�)v�.������+����y���iR��3���m�Ek�-@�傸��to�he�[���-� �,@��F�b"��j��e�F����̠��lv7�PZ� ��S�\Mӧ�aV��}��.Q�c�nV�����)�U�F����:̆w�i{��^�?	�=ӝ�<9A�M�F5O�[����~&���r�%��"*�T'�
��Iye��&fشĽ�z8��L�Z]�,�
��SڗG�S�kPW�����u0/�a��p��	���k�2��b�{�+T��(:�J��4�K	��Y46T�6V��g=��R�`�����a_�����ڡDI�I�8��K�����!��
G�RlDPq�2�'��`�~�G��H�ͬ��M���^휋���i	P��@�4��ܛdu{��/���O�i(PE>�RbDsM��Ʋ����}������G�Z԰[�\W_�"��֠���z�3[Ͻ�G��P���;qu*(��
�䱤��P�{%�'�g\�p����%��8����Ι���A�b���VH�-��5ݖS�V�N��)d a�s�0�8T��(<�D�;��._���vo���H��`aG ��إ��G�����NA�ޥp��58�}r��4�7�ڢA�?v#dCh�q�W����l����QKA���ֹ��l	��D���ז�~\�6���lW��q�PZ�|d�t'��Hb-F�z~�׍*_�v�#{1��z��%��j����!�!��D6��_n/��g���|I�# ��_j��{F{}E+�CGR��@�@u���EN�0c���M@ :R�is�z@���]j����X4<��K(8|�.b�)B9_�4�k2��83�_�.���� kг`	7���xU�z�&?�U�H[�s�=ųoA�Ef�t��F�,�)����2u�H����PU�Q�b���b�!�s�̭�꾭�>��._։
�9���(ȁ�{�,>S����+�1�~���͡@�����Hl�
!�����y�?�����`�
��ĳ��`ܷ-�8����HM�)=���K�����,|!��A�js:����x=!��3;�6=��T����|���dhJ���-�5���c �2��J4h]}$�u|�v� V�p3�杕 
�=L���뻁%p|�jƦ�����B֚��\��D?,�y����8Q�Q7��E��˵�e ѵ�����򭉅/}Rb��Yȴ�8so�z�.�E+>�1T2A�^3(�<����Z`Z�D>��a-$�wr� ��i������e})C��K���ߢ;�'Л��y�ck|��MbX�� )�e�J*�QA�z�*���BN +�wAP�j@3ߙSϓ<��/�G����qF�3���"짗-%�髩��^$+�.��)y+�
��b�:��a���h���]�M�3r����8/�9äLō	�X��/u� ��`���Ji��f��{.5d�	E9V����P:F5/T�K�Z�u�����۲���>}E�_E�� �ҝ5
��a�nZ�k��U?��kR򵾜4N��Q!�޸J茮�"Q�wր�!��1�$F^Y��!��>�G2/�ð��wy�+��j�1E9_��~D��d�FN@�<��n�'�/P[DQhH����S��K��F
fyY����-�����&{�@S�V��lcS"��.E��d���4�F�z�{���z �M�S�<���*m������.+�y�na��� �Rۉ�L����� Cu�f�g~��M7���������|.֐�
��$���(��)�Bu�!viLF:�ȡߩ�YJ�CQ;Px�İ�2~S�;���{Yx�m���T���O��Sk�T��\�ݳerU�Es���N��Zrг=-����+��Vְw���G�w70�(Tw�+�KX�{7�:�q�S�����w�A6�'y�O��0�	�G�7⛹[�.
�n��n�X�ɒ������mA�%�HH�@=�5����ݹ�$���"~��*�9 [��[4���=�VyR���Y�9�pK�� X������i����~^����$���@�0{����	�����q�_��ԐƧ��s�-Z�;ÑM� wl⼭�����/�/�Q�=MU�&� ����[W���K�� �� ��%�(z!>ɷvɾX�}�/=�(��OB�Ah)c�rdxM>f����>� ��A7�-�4����"
w���l;��H�	Ǔ�/�_�Q�i�b���+}�v��,�(M҄�+�ĪK��!X\���Bë�a�C�m���x������y���B
>����s�&���@���^�j0j�,��T��}�������H��-����_2;S����=&�NA��t����
V�G��q$�6Q�3r�=�HK�v	>L�k������I�t���\�{p�5���^i���&�ǖd	�D�-��=1w9�����S�+���RPzw�@k�Ãe�B�q�����'�tL��g�����/x��\B��;���S�	2���zӔㄓ#I�2󈣄��nԞWْ�^o�j�ɔ�gd݂j����]�&�O�����EDLo���s2[�kg6���w�%�-�t��C���e�{�%Ɗ��M_� ޒ�9|u��ޢm���߱���H
��'���ލđ��m���:�KEjJNz�=f��[�
��W�!�)� �-)�]�f�L���(���un��\-��������}k�l��mV7+f��Íu�~n��.Y<��,��Z�۵F �`�����ޔ�'0����� +5@�E�>�W֝I�{R��! J{���yo��0Yr��'�dzzvㅤ�!���a��p��f�!/ج�O�k�O<�U�W�	>�����g]�tZ�.ݝ�g_|�#A7�ń�b^X���Q]�/Z�.�3Y�m��%ˬc(�/�X×�m+~���s��j�`q@6&:Ґ��)���K��f#;�&�Wx��dh�?��YXA��f�2�ǶG���EW=��g��<��Np�	]��(P&���c���Er\��L����>�P"!;z�Nv�l�a�r�o���d~doʇ6�A�}<�c2��"�
�O9��`�ǀ��,�c�`y��IV���
���� \P|����jZ��5:\��~���]��8��=݈of@��s#��!�k��Q�w@��}��їw^�'�g�8c�"�����-`�g�y�ŧ�g�b���&'xWЋCQ}A�«i�/�CB��p�Hp&9�Y[<b�?���������֝��
,x!��H�xn�~�x���"ņ�¯{��=�v)vg�ٙ�љ�KjS3=��F$�7e9D�ho�w�^l��,A��V��5�������c��0�ǭN&���N��O���o� ����prd׷�R�b���I�e��s8Xh(ku��"�w�Y
7�9�8l ���Gl[��,��HgW_�ˡэq	?�L�6�@���,(hbl����4�Ж�B��y�dr
��O<Vۓ߉SQڈ�Q���):��ږ�)��V9�/���Rٍ�F���*Ff�[���@)_���q���GF�TK$@{���N������>�0�It@�WT%�Y���9�L��XlEB�ɱNW�Q]����_���+T��P$Ǡ^;�S}"%֘	"*ɇ���oS�2hP�7Q�� 6=7�g.|�uó�%���nk໘��7#�!��enNi�۾\�p��H,v<��b3��C�d�1��t)n쪆�+�,_��JD.�B�)��@ ����F7��60J��Be���>��L�2����|��j�Gھ��jp�v���Ɵ�53�dq�Q�sY
>{s�HWS���(���>���
rN6�I�H�=p��?�*�T��!��h=3��׻$I��%Z"�>�0D������褒���>��N��|�T�ؔ�^�Ϋ�F��K�b�c�&��Z+c⢲"�}�/ӵ�{�YD�]�`���dSК32�%D�ǐ�΍�!Nx���&����ET��p�	3�Z-�7���׉��^�������m�o�r�~
[b��6�W�Ď`���Se�%�m* ���oQ�/j��e�"zvv��Cz4	��),k�X��,`��Z,4�Gyc�c�bZ�sʌ�u8���s(�!'U����3�gY�khZ-ο���i�Fl[�Z��1�&�-��e��EE�>ӫ�o����?
.���=��5c���ZLl6�~�I�F���\�O��c&�cJ�uV�' ݘ���1�Y'm��>b�s�!,�MJ{.�~����I4��3��ClU�qW�<^�k�F����SH�|첝�5���]�v�����ZڞYYNaˈ�B=�Hfa�.�cT`܄k��|S]���g��4��0�C��	t]����r|E�n��e��Y��� �R�|w.�FOщ:�J���7��E���ت���Qhׁx(�N���V�H�����M&K�O��T^���9�- }�3$��E�3��I�Z��̦`�f���.&��.���4\��Z��^-��V�S���+7,(�K�r,@_z�Z���v�})�gVIL��͍�hu��q�S+�}OR�����9�Q�:g�pc44M�f�~wמe�x�)3� �G��w�-'�%�$k����u���~�w�k2J��v�#������QϛVa�R�q�(���Q�qH�]kW��C{����`��J�?o���V ظ�1�c�|��`������)�c����"�1��0*Ɠuo�
^Ԯ�\�{����ǁ>"�Gd����:�5o�C�%�� �v�ǜ:~���3'��a��.���;A!��:~Q]����\\^P�eIB�r���he�P�epo�������z�`$7ݡ'$EIu�4��v��_��*8���{�Q"�u:���[XW��>� T�����a13sN9���O��И9dO���r��tP����]�k->�0���J�}�
�P*j����s9Ѥ�l7��."�=�fDL����J谩3�^kU4�H��Ʊ�|�PtX�O`�I6��9�Iz��8�/��f�'u*Z��Yp��d�RC�١'���l!/�������{���0AP-Q�Ri<�$kl��ހʓD��=�?h�ݑx�&%[=����Hy�Ҩ/J���8�EC��{��-��;���,
B6�������J�sȻ��Ò�d�C����i���(b2�q�O�[��<�D�˹c�n���ЁG���Mi*r�'�hLG��|�F�oC����c5A4�o��Vf�}㝺�PǜX�l8�Xq���:�3��m�z�öQo���:g"D�:�v��W>�c����3� b�
�_�Y�-[ٍ�q&��@E�?&������1�Z�o ����R�." ����n`�.����Y̕ �Ԁh�z�|��ӯ�O�9�. (����1ݭ�D?�v�*�$��	�lT�?H�2T*���M��U��Sr��1x:L��C�"l��N	�Y�3դ�����n�Amh��	��=wyUqF�:}C�HV��#D�?�B<���A���KY�M�,�;�!��Z1uU������Q��K�8w�i(5��&f�_V*��� H�ֿ���2Gi�8��kfI���dk9tU1��nv3ĳ�@��.������Ng����k���^�!,� J:j=��V����t#�s՟�
K����D�1j�0p�}{=�R"�n��n�6	*	�5�<^����pN*]���7��C=\K�0�����H(�Z�*6!H+6����m���J]��m��Ө�LF/�O��.߀P�+�2=p�X�Y*��5�ɩ����Q"��Q�a�א(�Un���8���#���/��L�T��C<)��[(�Lֿ�-ȅ_kr0zi,	�=�a�B�tJ0�V�0���z�:�:}��������i�AgP�F ]v�'i�5]�[a	)�6!7EqN��1%�����eN9 �K%}��3肥2�1"�����snҦ�lI��Mz�@}��ލqr����}!p|��H�S�w�3r�#b��|m���7��.�����Y�����������p����@\|tT��2��ǻ4l��1��hqN򢦖d��sW����')�����Jo��.�nj��W�S���q����#b�3���.W�Л��9�$ٚ�%�K�X8�k=$j�j�y�n5COr�W�`JO�|öۊ��E�R�n}�$���Lֱ�zF�[����:@5��.}�Fd%�I0aZ+n��a�b�I͗(��&�16��d�*S:La��	uG��+��