��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���G�H�ƻ	�"�iQ�����3�7Q��㼫F|�ݽ0��@h ���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω��U��}��x�� �� ������[���a�8%`��4�s�6�XAoeu��a@����þ�V��1�Wqlw��9�K���m��+o���sp%��X�����b1Ø^���#K���lӧIA�a�V��R�5K�yQb�I����Gr�J�'�دv)h�V~�$v�p��"}�vo7k2a��pP.S��*����طǪh��p��U>?���>�`\��Yi���u����l�|���j@��"�O��$� ���xI+r�� 0�D�A�f�mXׂ�(ѳsv�`�S��Y�ix�P�Ra����+��a̞w���{ֱ@�W�8d4؇��2O��'HY-�z����s�1�WNcz7\F���r��RL�a))�kc�߇N	:.���n��{�'��?ɮ��N�7C��Hq-/��@�]\���<��9�`J�=�OLl??�L��y�����c��(r���U����i걲���9��m�!=�y����h�}y(;⟝*#rq��;nQ����>o?�M��;]/d^Bg�t��P	�x�[U���zy��<�hV�q��KPi8�����m��d�7������N\Q
7��0���Z�I��y�BR�J��?1;m�!=�y����h�}�Zn�h�>*��4D]�s�h6q3o?�M��;]��,��K!�ۻ2�e�1�ΟÈ�bHO���1���RL�a)r��fI���7+�.��sf���euw���wB"l��u���;��I�6r��f-Ӵv����N�Er��xXc)O�%�!�&��{G�3�^7����$������@���F���<r�O��C��0��`�R&.1��6��긲�7�M,0yV�u���;�j�g�v�*H�}����Ebzi`Ht����	x]�<���e��8�t�~��,�O�W��s�!5�S��H���)��������ҥ{E�?HF��eUٻo���mi��*	�ť�.^�i��' 1wH�x�xs��3�<A��z����
a�������~�+��,/,����W >g1�]l�&Y��F}갨y�����# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��`y��f2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�}�Z���ik2)�
}wʭU&H�1��8�h7H�u�ÍeRuw�C?3d,f$�7Q0�"<�F�ٴB�I�SbW�{b�2"���Bpш�#w��s8[Z�xZq��t�1�:�Ω�`<4}��o�r� ��J��ݪ��Ny5��	g�y�+��T��C�NJ���1�:�Ω�A��>s>;�t�  ",�r���q P�^�&d�A|�1�:�Ω��
�/�r�ѬL�1m��+5z�P�_X�I�?g�f�L#����2=�l�����4�c��ҁ����!��E���ƪϤ�Yk"1/��L�lW��+�va��2鍔�	g\A�Ny5��磋��w.V&��B֥�(����5�Z��f��Ո��D��2ER;�{m�B��,��B	hI�ˋ������Kp&�@���k�� ���3�ҺIÙ=�HgSmj�(����M���R��ӟ-��[7�d|���XP�����<��no#��٠R�^Ƒ���b9���j}8o{:��[MD|����a��'�-��띂ii�4];ˍH�P�(e�X�T}u��Q��L(\Ӧ�$�̎�)NC���)ҵ���]���>����C��ǩGY��-��%Mό���.ӳ�
�	?�<v�ј�"��Z鎬�������Ӊ*��y�7/����p���Z鎬����(��eظ���N:��e.��xu	���S8�/ #O�)R�^Ƒ����"X��[��Q[R�7�� ߌ�˕�(�
t��Y�{'%s���'����no#��٠R�^Ƒ����"X��[�'i�! ]���f�+��T�����h�6ؖ[!�� Q鹯e)�Op$!��o��R����r��X/��4�q�:�"��yȯS���Qߵs<��7�m��+e�(���n�JŬ+�"�却G�O��&�k��T:���V��9���Y��_E��V�no#��٠R�^Ƒ����"X��[��Q[R�7����n9�jsrCm�kO�=�ͦ�ڛ��4W�U����z~��6��	���`y����@����gG�[bGf�ޡ.pz�L�Y�{'%s���'����no#��٠R�^Ƒ����"X��[��&b2��sv��q͆c�!{p85��c���鿋�E~���W�6?��V���>?Mno#��٠R�^Ƒ��e>۵��>3R�d�ܦ)ݝOv%e�Vi���'�)�Բc��j*���F��
�D"�i:�gR���X��O���r����!�`�(i3����}��T��{���ʻ`�φ��<�6�@a� ���N����o�|�B��o��7�dPi��Y��bs��2[�a��o���Pi�#��R2W���R0s��>H�,b�z'hۉ)8D;�:㰻�߆�p�hؽ!�M��9�a>*<UB3 �~k�%�����Fodً���Fz�e<�Ia��la��o���Pi�#��Rq�\E��0谯n%�Z�'���Xw�j�7��+�uB;y��.U(�HN��R��#�mo�����Ě���R�`�)n�S߸��S�Ȍ`�*Ft���r%k$J&+��T�����D3���t�  ",�V��o5]�Q;�im��ȍry��	�
�I�>y!�`�(i3�І��%n3���bǆh�es��O��){�Ysy�t��P$u��&8�,�뼥<7.�G�p�P�hQ�GvEΡKCh��(	�G��^��AQ�0G�x#2���p[�Do�9�ҧ{�x����y�mZH֫&��5�q	�gh�䊉�䞘gx�n�W�����v;�k�@d���t��˳3[�u8�k/�z�xEQ���*[UxG�y��j��k
e�3+{�i�m�T�੉��%>�rG��M����{����"q�\E��0D������'���Xw�j�7��+�uB;y�Q[WG�i�D�wP�/�w,���^��5���ث	�+��r������@Z���rs�i���
(4��i�X���(㷾�N���H݆�